magic
tech sky130A
magscale 1 2
timestamp 1647565404
<< obsli1 >>
rect 1104 2159 73324 77265
<< obsm1 >>
rect 566 1572 73770 77296
<< metal2 >>
rect 1122 78800 1178 79600
rect 3422 78800 3478 79600
rect 5722 78800 5778 79600
rect 8022 78800 8078 79600
rect 10414 78800 10470 79600
rect 12714 78800 12770 79600
rect 15014 78800 15070 79600
rect 17314 78800 17370 79600
rect 19706 78800 19762 79600
rect 22006 78800 22062 79600
rect 24306 78800 24362 79600
rect 26698 78800 26754 79600
rect 28998 78800 29054 79600
rect 31298 78800 31354 79600
rect 33598 78800 33654 79600
rect 35990 78800 36046 79600
rect 38290 78800 38346 79600
rect 40590 78800 40646 79600
rect 42982 78800 43038 79600
rect 45282 78800 45338 79600
rect 47582 78800 47638 79600
rect 49882 78800 49938 79600
rect 52274 78800 52330 79600
rect 54574 78800 54630 79600
rect 56874 78800 56930 79600
rect 59266 78800 59322 79600
rect 61566 78800 61622 79600
rect 63866 78800 63922 79600
rect 66166 78800 66222 79600
rect 68558 78800 68614 79600
rect 70858 78800 70914 79600
rect 73158 78800 73214 79600
rect 570 0 626 800
rect 1766 0 1822 800
rect 2962 0 3018 800
rect 4158 0 4214 800
rect 5354 0 5410 800
rect 6550 0 6606 800
rect 7746 0 7802 800
rect 8942 0 8998 800
rect 10138 0 10194 800
rect 11334 0 11390 800
rect 12530 0 12586 800
rect 13726 0 13782 800
rect 14922 0 14978 800
rect 16118 0 16174 800
rect 17314 0 17370 800
rect 18510 0 18566 800
rect 19706 0 19762 800
rect 20902 0 20958 800
rect 22098 0 22154 800
rect 23294 0 23350 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 26974 0 27030 800
rect 28170 0 28226 800
rect 29366 0 29422 800
rect 30562 0 30618 800
rect 31758 0 31814 800
rect 32954 0 33010 800
rect 34150 0 34206 800
rect 35346 0 35402 800
rect 36542 0 36598 800
rect 37738 0 37794 800
rect 38934 0 38990 800
rect 40130 0 40186 800
rect 41326 0 41382 800
rect 42522 0 42578 800
rect 43718 0 43774 800
rect 44914 0 44970 800
rect 46110 0 46166 800
rect 47306 0 47362 800
rect 48502 0 48558 800
rect 49698 0 49754 800
rect 50986 0 51042 800
rect 52182 0 52238 800
rect 53378 0 53434 800
rect 54574 0 54630 800
rect 55770 0 55826 800
rect 56966 0 57022 800
rect 58162 0 58218 800
rect 59358 0 59414 800
rect 60554 0 60610 800
rect 61750 0 61806 800
rect 62946 0 63002 800
rect 64142 0 64198 800
rect 65338 0 65394 800
rect 66534 0 66590 800
rect 67730 0 67786 800
rect 68926 0 68982 800
rect 70122 0 70178 800
rect 71318 0 71374 800
rect 72514 0 72570 800
rect 73710 0 73766 800
<< obsm2 >>
rect 572 78744 1066 78962
rect 1234 78744 3366 78962
rect 3534 78744 5666 78962
rect 5834 78744 7966 78962
rect 8134 78744 10358 78962
rect 10526 78744 12658 78962
rect 12826 78744 14958 78962
rect 15126 78744 17258 78962
rect 17426 78744 19650 78962
rect 19818 78744 21950 78962
rect 22118 78744 24250 78962
rect 24418 78744 26642 78962
rect 26810 78744 28942 78962
rect 29110 78744 31242 78962
rect 31410 78744 33542 78962
rect 33710 78744 35934 78962
rect 36102 78744 38234 78962
rect 38402 78744 40534 78962
rect 40702 78744 42926 78962
rect 43094 78744 45226 78962
rect 45394 78744 47526 78962
rect 47694 78744 49826 78962
rect 49994 78744 52218 78962
rect 52386 78744 54518 78962
rect 54686 78744 56818 78962
rect 56986 78744 59210 78962
rect 59378 78744 61510 78962
rect 61678 78744 63810 78962
rect 63978 78744 66110 78962
rect 66278 78744 68502 78962
rect 68670 78744 70802 78962
rect 70970 78744 73102 78962
rect 73270 78744 73764 78962
rect 572 856 73764 78744
rect 682 575 1710 856
rect 1878 575 2906 856
rect 3074 575 4102 856
rect 4270 575 5298 856
rect 5466 575 6494 856
rect 6662 575 7690 856
rect 7858 575 8886 856
rect 9054 575 10082 856
rect 10250 575 11278 856
rect 11446 575 12474 856
rect 12642 575 13670 856
rect 13838 575 14866 856
rect 15034 575 16062 856
rect 16230 575 17258 856
rect 17426 575 18454 856
rect 18622 575 19650 856
rect 19818 575 20846 856
rect 21014 575 22042 856
rect 22210 575 23238 856
rect 23406 575 24434 856
rect 24602 575 25722 856
rect 25890 575 26918 856
rect 27086 575 28114 856
rect 28282 575 29310 856
rect 29478 575 30506 856
rect 30674 575 31702 856
rect 31870 575 32898 856
rect 33066 575 34094 856
rect 34262 575 35290 856
rect 35458 575 36486 856
rect 36654 575 37682 856
rect 37850 575 38878 856
rect 39046 575 40074 856
rect 40242 575 41270 856
rect 41438 575 42466 856
rect 42634 575 43662 856
rect 43830 575 44858 856
rect 45026 575 46054 856
rect 46222 575 47250 856
rect 47418 575 48446 856
rect 48614 575 49642 856
rect 49810 575 50930 856
rect 51098 575 52126 856
rect 52294 575 53322 856
rect 53490 575 54518 856
rect 54686 575 55714 856
rect 55882 575 56910 856
rect 57078 575 58106 856
rect 58274 575 59302 856
rect 59470 575 60498 856
rect 60666 575 61694 856
rect 61862 575 62890 856
rect 63058 575 64086 856
rect 64254 575 65282 856
rect 65450 575 66478 856
rect 66646 575 67674 856
rect 67842 575 68870 856
rect 69038 575 70066 856
rect 70234 575 71262 856
rect 71430 575 72458 856
rect 72626 575 73654 856
<< metal3 >>
rect 73670 78888 74470 79008
rect 0 78616 800 78736
rect 73670 77800 74470 77920
rect 0 76984 800 77104
rect 73670 76712 74470 76832
rect 73670 75624 74470 75744
rect 0 75216 800 75336
rect 73670 74400 74470 74520
rect 0 73584 800 73704
rect 73670 73312 74470 73432
rect 73670 72224 74470 72344
rect 0 71816 800 71936
rect 73670 71136 74470 71256
rect 0 70184 800 70304
rect 73670 69912 74470 70032
rect 73670 68824 74470 68944
rect 0 68416 800 68536
rect 73670 67736 74470 67856
rect 0 66784 800 66904
rect 73670 66648 74470 66768
rect 73670 65424 74470 65544
rect 0 65016 800 65136
rect 73670 64336 74470 64456
rect 0 63384 800 63504
rect 73670 63248 74470 63368
rect 73670 62160 74470 62280
rect 0 61752 800 61872
rect 73670 60936 74470 61056
rect 0 59984 800 60104
rect 73670 59848 74470 59968
rect 73670 58760 74470 58880
rect 0 58352 800 58472
rect 73670 57672 74470 57792
rect 0 56584 800 56704
rect 73670 56448 74470 56568
rect 73670 55360 74470 55480
rect 0 54952 800 55072
rect 73670 54272 74470 54392
rect 0 53184 800 53304
rect 73670 53184 74470 53304
rect 73670 52096 74470 52216
rect 0 51552 800 51672
rect 73670 50872 74470 50992
rect 0 49784 800 49904
rect 73670 49784 74470 49904
rect 73670 48696 74470 48816
rect 0 48152 800 48272
rect 73670 47608 74470 47728
rect 0 46520 800 46640
rect 73670 46384 74470 46504
rect 73670 45296 74470 45416
rect 0 44752 800 44872
rect 73670 44208 74470 44328
rect 0 43120 800 43240
rect 73670 43120 74470 43240
rect 73670 41896 74470 42016
rect 0 41352 800 41472
rect 73670 40808 74470 40928
rect 0 39720 800 39840
rect 73670 39720 74470 39840
rect 73670 38632 74470 38752
rect 0 37952 800 38072
rect 73670 37408 74470 37528
rect 0 36320 800 36440
rect 73670 36320 74470 36440
rect 73670 35232 74470 35352
rect 0 34552 800 34672
rect 73670 34144 74470 34264
rect 0 32920 800 33040
rect 73670 32920 74470 33040
rect 73670 31832 74470 31952
rect 0 31288 800 31408
rect 73670 30744 74470 30864
rect 0 29520 800 29640
rect 73670 29656 74470 29776
rect 73670 28432 74470 28552
rect 0 27888 800 28008
rect 73670 27344 74470 27464
rect 0 26120 800 26240
rect 73670 26256 74470 26376
rect 73670 25168 74470 25288
rect 0 24488 800 24608
rect 73670 24080 74470 24200
rect 0 22720 800 22840
rect 73670 22856 74470 22976
rect 73670 21768 74470 21888
rect 0 21088 800 21208
rect 73670 20680 74470 20800
rect 73670 19592 74470 19712
rect 0 19320 800 19440
rect 73670 18368 74470 18488
rect 0 17688 800 17808
rect 73670 17280 74470 17400
rect 0 16056 800 16176
rect 73670 16192 74470 16312
rect 73670 15104 74470 15224
rect 0 14288 800 14408
rect 73670 13880 74470 14000
rect 0 12656 800 12776
rect 73670 12792 74470 12912
rect 73670 11704 74470 11824
rect 0 10888 800 11008
rect 73670 10616 74470 10736
rect 0 9256 800 9376
rect 73670 9392 74470 9512
rect 73670 8304 74470 8424
rect 0 7488 800 7608
rect 73670 7216 74470 7336
rect 73670 6128 74470 6248
rect 0 5856 800 5976
rect 73670 4904 74470 5024
rect 0 4088 800 4208
rect 73670 3816 74470 3936
rect 73670 2728 74470 2848
rect 0 2456 800 2576
rect 73670 1640 74470 1760
rect 0 824 800 944
rect 73670 552 74470 672
<< obsm3 >>
rect 800 77184 73670 77281
rect 880 76912 73670 77184
rect 880 76904 73590 76912
rect 800 76632 73590 76904
rect 800 75824 73670 76632
rect 800 75544 73590 75824
rect 800 75416 73670 75544
rect 880 75136 73670 75416
rect 800 74600 73670 75136
rect 800 74320 73590 74600
rect 800 73784 73670 74320
rect 880 73512 73670 73784
rect 880 73504 73590 73512
rect 800 73232 73590 73504
rect 800 72424 73670 73232
rect 800 72144 73590 72424
rect 800 72016 73670 72144
rect 880 71736 73670 72016
rect 800 71336 73670 71736
rect 800 71056 73590 71336
rect 800 70384 73670 71056
rect 880 70112 73670 70384
rect 880 70104 73590 70112
rect 800 69832 73590 70104
rect 800 69024 73670 69832
rect 800 68744 73590 69024
rect 800 68616 73670 68744
rect 880 68336 73670 68616
rect 800 67936 73670 68336
rect 800 67656 73590 67936
rect 800 66984 73670 67656
rect 880 66848 73670 66984
rect 880 66704 73590 66848
rect 800 66568 73590 66704
rect 800 65624 73670 66568
rect 800 65344 73590 65624
rect 800 65216 73670 65344
rect 880 64936 73670 65216
rect 800 64536 73670 64936
rect 800 64256 73590 64536
rect 800 63584 73670 64256
rect 880 63448 73670 63584
rect 880 63304 73590 63448
rect 800 63168 73590 63304
rect 800 62360 73670 63168
rect 800 62080 73590 62360
rect 800 61952 73670 62080
rect 880 61672 73670 61952
rect 800 61136 73670 61672
rect 800 60856 73590 61136
rect 800 60184 73670 60856
rect 880 60048 73670 60184
rect 880 59904 73590 60048
rect 800 59768 73590 59904
rect 800 58960 73670 59768
rect 800 58680 73590 58960
rect 800 58552 73670 58680
rect 880 58272 73670 58552
rect 800 57872 73670 58272
rect 800 57592 73590 57872
rect 800 56784 73670 57592
rect 880 56648 73670 56784
rect 880 56504 73590 56648
rect 800 56368 73590 56504
rect 800 55560 73670 56368
rect 800 55280 73590 55560
rect 800 55152 73670 55280
rect 880 54872 73670 55152
rect 800 54472 73670 54872
rect 800 54192 73590 54472
rect 800 53384 73670 54192
rect 880 53104 73590 53384
rect 800 52296 73670 53104
rect 800 52016 73590 52296
rect 800 51752 73670 52016
rect 880 51472 73670 51752
rect 800 51072 73670 51472
rect 800 50792 73590 51072
rect 800 49984 73670 50792
rect 880 49704 73590 49984
rect 800 48896 73670 49704
rect 800 48616 73590 48896
rect 800 48352 73670 48616
rect 880 48072 73670 48352
rect 800 47808 73670 48072
rect 800 47528 73590 47808
rect 800 46720 73670 47528
rect 880 46584 73670 46720
rect 880 46440 73590 46584
rect 800 46304 73590 46440
rect 800 45496 73670 46304
rect 800 45216 73590 45496
rect 800 44952 73670 45216
rect 880 44672 73670 44952
rect 800 44408 73670 44672
rect 800 44128 73590 44408
rect 800 43320 73670 44128
rect 880 43040 73590 43320
rect 800 42096 73670 43040
rect 800 41816 73590 42096
rect 800 41552 73670 41816
rect 880 41272 73670 41552
rect 800 41008 73670 41272
rect 800 40728 73590 41008
rect 800 39920 73670 40728
rect 880 39640 73590 39920
rect 800 38832 73670 39640
rect 800 38552 73590 38832
rect 800 38152 73670 38552
rect 880 37872 73670 38152
rect 800 37608 73670 37872
rect 800 37328 73590 37608
rect 800 36520 73670 37328
rect 880 36240 73590 36520
rect 800 35432 73670 36240
rect 800 35152 73590 35432
rect 800 34752 73670 35152
rect 880 34472 73670 34752
rect 800 34344 73670 34472
rect 800 34064 73590 34344
rect 800 33120 73670 34064
rect 880 32840 73590 33120
rect 800 32032 73670 32840
rect 800 31752 73590 32032
rect 800 31488 73670 31752
rect 880 31208 73670 31488
rect 800 30944 73670 31208
rect 800 30664 73590 30944
rect 800 29856 73670 30664
rect 800 29720 73590 29856
rect 880 29576 73590 29720
rect 880 29440 73670 29576
rect 800 28632 73670 29440
rect 800 28352 73590 28632
rect 800 28088 73670 28352
rect 880 27808 73670 28088
rect 800 27544 73670 27808
rect 800 27264 73590 27544
rect 800 26456 73670 27264
rect 800 26320 73590 26456
rect 880 26176 73590 26320
rect 880 26040 73670 26176
rect 800 25368 73670 26040
rect 800 25088 73590 25368
rect 800 24688 73670 25088
rect 880 24408 73670 24688
rect 800 24280 73670 24408
rect 800 24000 73590 24280
rect 800 23056 73670 24000
rect 800 22920 73590 23056
rect 880 22776 73590 22920
rect 880 22640 73670 22776
rect 800 21968 73670 22640
rect 800 21688 73590 21968
rect 800 21288 73670 21688
rect 880 21008 73670 21288
rect 800 20880 73670 21008
rect 800 20600 73590 20880
rect 800 19792 73670 20600
rect 800 19520 73590 19792
rect 880 19512 73590 19520
rect 880 19240 73670 19512
rect 800 18568 73670 19240
rect 800 18288 73590 18568
rect 800 17888 73670 18288
rect 880 17608 73670 17888
rect 800 17480 73670 17608
rect 800 17200 73590 17480
rect 800 16392 73670 17200
rect 800 16256 73590 16392
rect 880 16112 73590 16256
rect 880 15976 73670 16112
rect 800 15304 73670 15976
rect 800 15024 73590 15304
rect 800 14488 73670 15024
rect 880 14208 73670 14488
rect 800 14080 73670 14208
rect 800 13800 73590 14080
rect 800 12992 73670 13800
rect 800 12856 73590 12992
rect 880 12712 73590 12856
rect 880 12576 73670 12712
rect 800 11904 73670 12576
rect 800 11624 73590 11904
rect 800 11088 73670 11624
rect 880 10816 73670 11088
rect 880 10808 73590 10816
rect 800 10536 73590 10808
rect 800 9592 73670 10536
rect 800 9456 73590 9592
rect 880 9312 73590 9456
rect 880 9176 73670 9312
rect 800 8504 73670 9176
rect 800 8224 73590 8504
rect 800 7688 73670 8224
rect 880 7416 73670 7688
rect 880 7408 73590 7416
rect 800 7136 73590 7408
rect 800 6328 73670 7136
rect 800 6056 73590 6328
rect 880 6048 73590 6056
rect 880 5776 73670 6048
rect 800 5104 73670 5776
rect 800 4824 73590 5104
rect 800 4288 73670 4824
rect 880 4016 73670 4288
rect 880 4008 73590 4016
rect 800 3736 73590 4008
rect 800 2928 73670 3736
rect 800 2656 73590 2928
rect 880 2648 73590 2656
rect 880 2376 73670 2648
rect 800 1840 73670 2376
rect 800 1560 73590 1840
rect 800 1024 73670 1560
rect 880 752 73670 1024
rect 880 744 73590 752
rect 800 579 73590 744
<< metal4 >>
rect 4208 2128 4528 77296
rect 19568 2128 19888 77296
rect 34928 2128 35248 77296
rect 50288 2128 50608 77296
rect 65648 2128 65968 77296
<< obsm4 >>
rect 2083 3027 4128 76941
rect 4608 3027 19488 76941
rect 19968 3027 34848 76941
rect 35328 3027 50208 76941
rect 50688 3027 65568 76941
rect 66048 3027 71517 76941
<< labels >>
rlabel metal2 s 570 0 626 800 6 active
port 1 nsew signal input
rlabel metal3 s 73670 67736 74470 67856 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 12714 78800 12770 79600 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 10414 78800 10470 79600 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 8022 78800 8078 79600 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 5722 78800 5778 79600 6 io_in[13]
port 6 nsew signal input
rlabel metal3 s 73670 56448 74470 56568 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 73670 55360 74470 55480 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 3422 78800 3478 79600 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 1122 78800 1178 79600 6 io_in[17]
port 10 nsew signal input
rlabel metal3 s 73670 11704 74470 11824 6 io_in[18]
port 11 nsew signal input
rlabel metal3 s 73670 10616 74470 10736 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 73670 66648 74470 66768 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 73670 54272 74470 54392 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 73670 53184 74470 53304 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 73670 9392 74470 9512 6 io_in[22]
port 16 nsew signal input
rlabel metal3 s 73670 8304 74470 8424 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 73670 7216 74470 7336 6 io_in[24]
port 18 nsew signal input
rlabel metal3 s 73670 6128 74470 6248 6 io_in[25]
port 19 nsew signal input
rlabel metal3 s 73670 4904 74470 5024 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 73670 52096 74470 52216 6 io_in[27]
port 21 nsew signal input
rlabel metal3 s 73670 50872 74470 50992 6 io_in[28]
port 22 nsew signal input
rlabel metal3 s 73670 49784 74470 49904 6 io_in[29]
port 23 nsew signal input
rlabel metal3 s 73670 65424 74470 65544 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 73670 3816 74470 3936 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 73670 2728 74470 2848 6 io_in[31]
port 26 nsew signal input
rlabel metal3 s 73670 1640 74470 1760 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 73670 552 74470 672 6 io_in[33]
port 28 nsew signal input
rlabel metal3 s 73670 48696 74470 48816 6 io_in[34]
port 29 nsew signal input
rlabel metal3 s 73670 47608 74470 47728 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 73670 46384 74470 46504 6 io_in[36]
port 31 nsew signal input
rlabel metal3 s 73670 45296 74470 45416 6 io_in[37]
port 32 nsew signal input
rlabel metal3 s 73670 64336 74470 64456 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 73670 63248 74470 63368 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 73670 62160 74470 62280 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 73670 60936 74470 61056 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 73670 59848 74470 59968 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 73670 58760 74470 58880 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 73670 57672 74470 57792 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 io_oeb[16]
port 47 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 io_oeb[17]
port 48 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 0 824 800 944 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 73158 78800 73214 79600 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 70858 78800 70914 79600 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 68558 78800 68614 79600 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 66166 78800 66222 79600 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 63866 78800 63922 79600 6 io_oeb[25]
port 57 nsew signal output
rlabel metal2 s 61566 78800 61622 79600 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 59266 78800 59322 79600 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 56874 78800 56930 79600 6 io_oeb[28]
port 60 nsew signal output
rlabel metal2 s 54574 78800 54630 79600 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 52274 78800 52330 79600 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 49882 78800 49938 79600 6 io_oeb[31]
port 64 nsew signal output
rlabel metal2 s 47582 78800 47638 79600 6 io_oeb[32]
port 65 nsew signal output
rlabel metal2 s 45282 78800 45338 79600 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 42982 78800 43038 79600 6 io_oeb[34]
port 67 nsew signal output
rlabel metal2 s 40590 78800 40646 79600 6 io_oeb[35]
port 68 nsew signal output
rlabel metal2 s 38290 78800 38346 79600 6 io_oeb[36]
port 69 nsew signal output
rlabel metal2 s 35990 78800 36046 79600 6 io_oeb[37]
port 70 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 73670 44208 74470 44328 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 73670 32920 74470 33040 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 73670 31832 74470 31952 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 73670 30744 74470 30864 6 io_out[12]
port 81 nsew signal output
rlabel metal3 s 73670 29656 74470 29776 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 73670 28432 74470 28552 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 73670 27344 74470 27464 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 73670 26256 74470 26376 6 io_out[16]
port 85 nsew signal output
rlabel metal3 s 73670 25168 74470 25288 6 io_out[17]
port 86 nsew signal output
rlabel metal3 s 73670 24080 74470 24200 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 73670 22856 74470 22976 6 io_out[19]
port 88 nsew signal output
rlabel metal3 s 73670 43120 74470 43240 6 io_out[1]
port 89 nsew signal output
rlabel metal3 s 73670 21768 74470 21888 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 73670 20680 74470 20800 6 io_out[21]
port 91 nsew signal output
rlabel metal3 s 73670 19592 74470 19712 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 73670 18368 74470 18488 6 io_out[23]
port 93 nsew signal output
rlabel metal3 s 73670 17280 74470 17400 6 io_out[24]
port 94 nsew signal output
rlabel metal3 s 73670 16192 74470 16312 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 73670 15104 74470 15224 6 io_out[26]
port 96 nsew signal output
rlabel metal3 s 73670 13880 74470 14000 6 io_out[27]
port 97 nsew signal output
rlabel metal3 s 73670 12792 74470 12912 6 io_out[28]
port 98 nsew signal output
rlabel metal2 s 33598 78800 33654 79600 6 io_out[29]
port 99 nsew signal output
rlabel metal3 s 73670 41896 74470 42016 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 31298 78800 31354 79600 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 28998 78800 29054 79600 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 26698 78800 26754 79600 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 24306 78800 24362 79600 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 22006 78800 22062 79600 6 io_out[34]
port 105 nsew signal output
rlabel metal2 s 19706 78800 19762 79600 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 17314 78800 17370 79600 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 15014 78800 15070 79600 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 73670 40808 74470 40928 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 73670 39720 74470 39840 6 io_out[4]
port 110 nsew signal output
rlabel metal3 s 73670 38632 74470 38752 6 io_out[5]
port 111 nsew signal output
rlabel metal3 s 73670 37408 74470 37528 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 73670 36320 74470 36440 6 io_out[7]
port 113 nsew signal output
rlabel metal3 s 73670 35232 74470 35352 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 73670 34144 74470 34264 6 io_out[9]
port 115 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 73670 72224 74470 72344 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 73670 71136 74470 71256 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 73670 69912 74470 70032 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 73670 68824 74470 68944 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal2 s 59358 0 59414 800 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal2 s 42522 0 42578 800 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal2 s 66534 0 66590 800 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 0 59984 800 60104 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal3 s 0 53184 800 53304 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 73670 78888 74470 79008 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 73670 77800 74470 77920 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 73670 76712 74470 76832 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 73670 75624 74470 75744 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 73670 74400 74470 74520 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 73670 73312 74470 73432 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 2128 4528 77296 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 2128 35248 77296 6 vccd1
port 212 nsew power input
rlabel metal4 s 65648 2128 65968 77296 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 2128 19888 77296 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 2128 50608 77296 6 vssd1
port 213 nsew ground input
rlabel metal2 s 1766 0 1822 800 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 74470 79600
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 17379296
string GDS_FILE /openlane/designs/wrapped_hack_soc_dffram/runs/RUN_2022.03.18_00.58.38/results/finishing/wrapped_hack_soc_dffram.magic.gds
string GDS_START 9615550
<< end >>

