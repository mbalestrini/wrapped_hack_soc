magic
tech sky130A
magscale 1 2
timestamp 1647447067
<< obsli1 >>
rect 989 2159 77280 77265
<< obsm1 >>
rect 566 1708 77818 77296
<< metal2 >>
rect 1214 78800 1270 79600
rect 3606 78800 3662 79600
rect 6090 78800 6146 79600
rect 8482 78800 8538 79600
rect 10966 78800 11022 79600
rect 13450 78800 13506 79600
rect 15842 78800 15898 79600
rect 18326 78800 18382 79600
rect 20810 78800 20866 79600
rect 23202 78800 23258 79600
rect 25686 78800 25742 79600
rect 28170 78800 28226 79600
rect 30562 78800 30618 79600
rect 33046 78800 33102 79600
rect 35530 78800 35586 79600
rect 37922 78800 37978 79600
rect 40406 78800 40462 79600
rect 42890 78800 42946 79600
rect 45282 78800 45338 79600
rect 47766 78800 47822 79600
rect 50250 78800 50306 79600
rect 52642 78800 52698 79600
rect 55126 78800 55182 79600
rect 57610 78800 57666 79600
rect 60002 78800 60058 79600
rect 62486 78800 62542 79600
rect 64970 78800 65026 79600
rect 67362 78800 67418 79600
rect 69846 78800 69902 79600
rect 72330 78800 72386 79600
rect 74722 78800 74778 79600
rect 77206 78800 77262 79600
rect 570 0 626 800
rect 1766 0 1822 800
rect 3054 0 3110 800
rect 4342 0 4398 800
rect 5630 0 5686 800
rect 6826 0 6882 800
rect 8114 0 8170 800
rect 9402 0 9458 800
rect 10690 0 10746 800
rect 11886 0 11942 800
rect 13174 0 13230 800
rect 14462 0 14518 800
rect 15750 0 15806 800
rect 16946 0 17002 800
rect 18234 0 18290 800
rect 19522 0 19578 800
rect 20810 0 20866 800
rect 22006 0 22062 800
rect 23294 0 23350 800
rect 24582 0 24638 800
rect 25870 0 25926 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 30930 0 30986 800
rect 32126 0 32182 800
rect 33414 0 33470 800
rect 34702 0 34758 800
rect 35990 0 36046 800
rect 37186 0 37242 800
rect 38474 0 38530 800
rect 39762 0 39818 800
rect 41050 0 41106 800
rect 42338 0 42394 800
rect 43534 0 43590 800
rect 44822 0 44878 800
rect 46110 0 46166 800
rect 47398 0 47454 800
rect 48594 0 48650 800
rect 49882 0 49938 800
rect 51170 0 51226 800
rect 52458 0 52514 800
rect 53654 0 53710 800
rect 54942 0 54998 800
rect 56230 0 56286 800
rect 57518 0 57574 800
rect 58714 0 58770 800
rect 60002 0 60058 800
rect 61290 0 61346 800
rect 62578 0 62634 800
rect 63774 0 63830 800
rect 65062 0 65118 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68834 0 68890 800
rect 70122 0 70178 800
rect 71410 0 71466 800
rect 72698 0 72754 800
rect 73894 0 73950 800
rect 75182 0 75238 800
rect 76470 0 76526 800
rect 77758 0 77814 800
<< obsm2 >>
rect 572 78744 1158 78962
rect 1326 78744 3550 78962
rect 3718 78744 6034 78962
rect 6202 78744 8426 78962
rect 8594 78744 10910 78962
rect 11078 78744 13394 78962
rect 13562 78744 15786 78962
rect 15954 78744 18270 78962
rect 18438 78744 20754 78962
rect 20922 78744 23146 78962
rect 23314 78744 25630 78962
rect 25798 78744 28114 78962
rect 28282 78744 30506 78962
rect 30674 78744 32990 78962
rect 33158 78744 35474 78962
rect 35642 78744 37866 78962
rect 38034 78744 40350 78962
rect 40518 78744 42834 78962
rect 43002 78744 45226 78962
rect 45394 78744 47710 78962
rect 47878 78744 50194 78962
rect 50362 78744 52586 78962
rect 52754 78744 55070 78962
rect 55238 78744 57554 78962
rect 57722 78744 59946 78962
rect 60114 78744 62430 78962
rect 62598 78744 64914 78962
rect 65082 78744 67306 78962
rect 67474 78744 69790 78962
rect 69958 78744 72274 78962
rect 72442 78744 74666 78962
rect 74834 78744 77150 78962
rect 77318 78744 77812 78962
rect 572 856 77812 78744
rect 682 575 1710 856
rect 1878 575 2998 856
rect 3166 575 4286 856
rect 4454 575 5574 856
rect 5742 575 6770 856
rect 6938 575 8058 856
rect 8226 575 9346 856
rect 9514 575 10634 856
rect 10802 575 11830 856
rect 11998 575 13118 856
rect 13286 575 14406 856
rect 14574 575 15694 856
rect 15862 575 16890 856
rect 17058 575 18178 856
rect 18346 575 19466 856
rect 19634 575 20754 856
rect 20922 575 21950 856
rect 22118 575 23238 856
rect 23406 575 24526 856
rect 24694 575 25814 856
rect 25982 575 27010 856
rect 27178 575 28298 856
rect 28466 575 29586 856
rect 29754 575 30874 856
rect 31042 575 32070 856
rect 32238 575 33358 856
rect 33526 575 34646 856
rect 34814 575 35934 856
rect 36102 575 37130 856
rect 37298 575 38418 856
rect 38586 575 39706 856
rect 39874 575 40994 856
rect 41162 575 42282 856
rect 42450 575 43478 856
rect 43646 575 44766 856
rect 44934 575 46054 856
rect 46222 575 47342 856
rect 47510 575 48538 856
rect 48706 575 49826 856
rect 49994 575 51114 856
rect 51282 575 52402 856
rect 52570 575 53598 856
rect 53766 575 54886 856
rect 55054 575 56174 856
rect 56342 575 57462 856
rect 57630 575 58658 856
rect 58826 575 59946 856
rect 60114 575 61234 856
rect 61402 575 62522 856
rect 62690 575 63718 856
rect 63886 575 65006 856
rect 65174 575 66294 856
rect 66462 575 67582 856
rect 67750 575 68778 856
rect 68946 575 70066 856
rect 70234 575 71354 856
rect 71522 575 72642 856
rect 72810 575 73838 856
rect 74006 575 75126 856
rect 75294 575 76414 856
rect 76582 575 77702 856
<< metal3 >>
rect 77650 78888 78450 79008
rect 0 78616 800 78736
rect 77650 77800 78450 77920
rect 0 76984 800 77104
rect 77650 76712 78450 76832
rect 77650 75624 78450 75744
rect 0 75216 800 75336
rect 77650 74400 78450 74520
rect 0 73584 800 73704
rect 77650 73312 78450 73432
rect 77650 72224 78450 72344
rect 0 71816 800 71936
rect 77650 71136 78450 71256
rect 0 70184 800 70304
rect 77650 69912 78450 70032
rect 77650 68824 78450 68944
rect 0 68416 800 68536
rect 77650 67736 78450 67856
rect 0 66784 800 66904
rect 77650 66648 78450 66768
rect 77650 65424 78450 65544
rect 0 65016 800 65136
rect 77650 64336 78450 64456
rect 0 63384 800 63504
rect 77650 63248 78450 63368
rect 77650 62160 78450 62280
rect 0 61752 800 61872
rect 77650 60936 78450 61056
rect 0 59984 800 60104
rect 77650 59848 78450 59968
rect 77650 58760 78450 58880
rect 0 58352 800 58472
rect 77650 57672 78450 57792
rect 0 56584 800 56704
rect 77650 56448 78450 56568
rect 77650 55360 78450 55480
rect 0 54952 800 55072
rect 77650 54272 78450 54392
rect 0 53184 800 53304
rect 77650 53184 78450 53304
rect 77650 52096 78450 52216
rect 0 51552 800 51672
rect 77650 50872 78450 50992
rect 0 49784 800 49904
rect 77650 49784 78450 49904
rect 77650 48696 78450 48816
rect 0 48152 800 48272
rect 77650 47608 78450 47728
rect 0 46520 800 46640
rect 77650 46384 78450 46504
rect 77650 45296 78450 45416
rect 0 44752 800 44872
rect 77650 44208 78450 44328
rect 0 43120 800 43240
rect 77650 43120 78450 43240
rect 77650 41896 78450 42016
rect 0 41352 800 41472
rect 77650 40808 78450 40928
rect 0 39720 800 39840
rect 77650 39720 78450 39840
rect 77650 38632 78450 38752
rect 0 37952 800 38072
rect 77650 37408 78450 37528
rect 0 36320 800 36440
rect 77650 36320 78450 36440
rect 77650 35232 78450 35352
rect 0 34552 800 34672
rect 77650 34144 78450 34264
rect 0 32920 800 33040
rect 77650 32920 78450 33040
rect 77650 31832 78450 31952
rect 0 31288 800 31408
rect 77650 30744 78450 30864
rect 0 29520 800 29640
rect 77650 29656 78450 29776
rect 77650 28432 78450 28552
rect 0 27888 800 28008
rect 77650 27344 78450 27464
rect 0 26120 800 26240
rect 77650 26256 78450 26376
rect 77650 25168 78450 25288
rect 0 24488 800 24608
rect 77650 24080 78450 24200
rect 0 22720 800 22840
rect 77650 22856 78450 22976
rect 77650 21768 78450 21888
rect 0 21088 800 21208
rect 77650 20680 78450 20800
rect 77650 19592 78450 19712
rect 0 19320 800 19440
rect 77650 18368 78450 18488
rect 0 17688 800 17808
rect 77650 17280 78450 17400
rect 0 16056 800 16176
rect 77650 16192 78450 16312
rect 77650 15104 78450 15224
rect 0 14288 800 14408
rect 77650 13880 78450 14000
rect 0 12656 800 12776
rect 77650 12792 78450 12912
rect 77650 11704 78450 11824
rect 0 10888 800 11008
rect 77650 10616 78450 10736
rect 0 9256 800 9376
rect 77650 9392 78450 9512
rect 77650 8304 78450 8424
rect 0 7488 800 7608
rect 77650 7216 78450 7336
rect 77650 6128 78450 6248
rect 0 5856 800 5976
rect 77650 4904 78450 5024
rect 0 4088 800 4208
rect 77650 3816 78450 3936
rect 77650 2728 78450 2848
rect 0 2456 800 2576
rect 77650 1640 78450 1760
rect 0 824 800 944
rect 77650 552 78450 672
<< obsm3 >>
rect 800 77184 77650 77281
rect 880 76912 77650 77184
rect 880 76904 77570 76912
rect 800 76632 77570 76904
rect 800 75824 77650 76632
rect 800 75544 77570 75824
rect 800 75416 77650 75544
rect 880 75136 77650 75416
rect 800 74600 77650 75136
rect 800 74320 77570 74600
rect 800 73784 77650 74320
rect 880 73512 77650 73784
rect 880 73504 77570 73512
rect 800 73232 77570 73504
rect 800 72424 77650 73232
rect 800 72144 77570 72424
rect 800 72016 77650 72144
rect 880 71736 77650 72016
rect 800 71336 77650 71736
rect 800 71056 77570 71336
rect 800 70384 77650 71056
rect 880 70112 77650 70384
rect 880 70104 77570 70112
rect 800 69832 77570 70104
rect 800 69024 77650 69832
rect 800 68744 77570 69024
rect 800 68616 77650 68744
rect 880 68336 77650 68616
rect 800 67936 77650 68336
rect 800 67656 77570 67936
rect 800 66984 77650 67656
rect 880 66848 77650 66984
rect 880 66704 77570 66848
rect 800 66568 77570 66704
rect 800 65624 77650 66568
rect 800 65344 77570 65624
rect 800 65216 77650 65344
rect 880 64936 77650 65216
rect 800 64536 77650 64936
rect 800 64256 77570 64536
rect 800 63584 77650 64256
rect 880 63448 77650 63584
rect 880 63304 77570 63448
rect 800 63168 77570 63304
rect 800 62360 77650 63168
rect 800 62080 77570 62360
rect 800 61952 77650 62080
rect 880 61672 77650 61952
rect 800 61136 77650 61672
rect 800 60856 77570 61136
rect 800 60184 77650 60856
rect 880 60048 77650 60184
rect 880 59904 77570 60048
rect 800 59768 77570 59904
rect 800 58960 77650 59768
rect 800 58680 77570 58960
rect 800 58552 77650 58680
rect 880 58272 77650 58552
rect 800 57872 77650 58272
rect 800 57592 77570 57872
rect 800 56784 77650 57592
rect 880 56648 77650 56784
rect 880 56504 77570 56648
rect 800 56368 77570 56504
rect 800 55560 77650 56368
rect 800 55280 77570 55560
rect 800 55152 77650 55280
rect 880 54872 77650 55152
rect 800 54472 77650 54872
rect 800 54192 77570 54472
rect 800 53384 77650 54192
rect 880 53104 77570 53384
rect 800 52296 77650 53104
rect 800 52016 77570 52296
rect 800 51752 77650 52016
rect 880 51472 77650 51752
rect 800 51072 77650 51472
rect 800 50792 77570 51072
rect 800 49984 77650 50792
rect 880 49704 77570 49984
rect 800 48896 77650 49704
rect 800 48616 77570 48896
rect 800 48352 77650 48616
rect 880 48072 77650 48352
rect 800 47808 77650 48072
rect 800 47528 77570 47808
rect 800 46720 77650 47528
rect 880 46584 77650 46720
rect 880 46440 77570 46584
rect 800 46304 77570 46440
rect 800 45496 77650 46304
rect 800 45216 77570 45496
rect 800 44952 77650 45216
rect 880 44672 77650 44952
rect 800 44408 77650 44672
rect 800 44128 77570 44408
rect 800 43320 77650 44128
rect 880 43040 77570 43320
rect 800 42096 77650 43040
rect 800 41816 77570 42096
rect 800 41552 77650 41816
rect 880 41272 77650 41552
rect 800 41008 77650 41272
rect 800 40728 77570 41008
rect 800 39920 77650 40728
rect 880 39640 77570 39920
rect 800 38832 77650 39640
rect 800 38552 77570 38832
rect 800 38152 77650 38552
rect 880 37872 77650 38152
rect 800 37608 77650 37872
rect 800 37328 77570 37608
rect 800 36520 77650 37328
rect 880 36240 77570 36520
rect 800 35432 77650 36240
rect 800 35152 77570 35432
rect 800 34752 77650 35152
rect 880 34472 77650 34752
rect 800 34344 77650 34472
rect 800 34064 77570 34344
rect 800 33120 77650 34064
rect 880 32840 77570 33120
rect 800 32032 77650 32840
rect 800 31752 77570 32032
rect 800 31488 77650 31752
rect 880 31208 77650 31488
rect 800 30944 77650 31208
rect 800 30664 77570 30944
rect 800 29856 77650 30664
rect 800 29720 77570 29856
rect 880 29576 77570 29720
rect 880 29440 77650 29576
rect 800 28632 77650 29440
rect 800 28352 77570 28632
rect 800 28088 77650 28352
rect 880 27808 77650 28088
rect 800 27544 77650 27808
rect 800 27264 77570 27544
rect 800 26456 77650 27264
rect 800 26320 77570 26456
rect 880 26176 77570 26320
rect 880 26040 77650 26176
rect 800 25368 77650 26040
rect 800 25088 77570 25368
rect 800 24688 77650 25088
rect 880 24408 77650 24688
rect 800 24280 77650 24408
rect 800 24000 77570 24280
rect 800 23056 77650 24000
rect 800 22920 77570 23056
rect 880 22776 77570 22920
rect 880 22640 77650 22776
rect 800 21968 77650 22640
rect 800 21688 77570 21968
rect 800 21288 77650 21688
rect 880 21008 77650 21288
rect 800 20880 77650 21008
rect 800 20600 77570 20880
rect 800 19792 77650 20600
rect 800 19520 77570 19792
rect 880 19512 77570 19520
rect 880 19240 77650 19512
rect 800 18568 77650 19240
rect 800 18288 77570 18568
rect 800 17888 77650 18288
rect 880 17608 77650 17888
rect 800 17480 77650 17608
rect 800 17200 77570 17480
rect 800 16392 77650 17200
rect 800 16256 77570 16392
rect 880 16112 77570 16256
rect 880 15976 77650 16112
rect 800 15304 77650 15976
rect 800 15024 77570 15304
rect 800 14488 77650 15024
rect 880 14208 77650 14488
rect 800 14080 77650 14208
rect 800 13800 77570 14080
rect 800 12992 77650 13800
rect 800 12856 77570 12992
rect 880 12712 77570 12856
rect 880 12576 77650 12712
rect 800 11904 77650 12576
rect 800 11624 77570 11904
rect 800 11088 77650 11624
rect 880 10816 77650 11088
rect 880 10808 77570 10816
rect 800 10536 77570 10808
rect 800 9592 77650 10536
rect 800 9456 77570 9592
rect 880 9312 77570 9456
rect 880 9176 77650 9312
rect 800 8504 77650 9176
rect 800 8224 77570 8504
rect 800 7688 77650 8224
rect 880 7416 77650 7688
rect 880 7408 77570 7416
rect 800 7136 77570 7408
rect 800 6328 77650 7136
rect 800 6056 77570 6328
rect 880 6048 77570 6056
rect 880 5776 77650 6048
rect 800 5104 77650 5776
rect 800 4824 77570 5104
rect 800 4288 77650 4824
rect 880 4016 77650 4288
rect 880 4008 77570 4016
rect 800 3736 77570 4008
rect 800 2928 77650 3736
rect 800 2656 77570 2928
rect 880 2648 77570 2656
rect 880 2376 77650 2648
rect 800 1840 77650 2376
rect 800 1560 77570 1840
rect 800 1024 77650 1560
rect 880 752 77650 1024
rect 880 744 77570 752
rect 800 579 77570 744
<< metal4 >>
rect 4208 2128 4528 77296
rect 19568 2128 19888 77296
rect 34928 2128 35248 77296
rect 50288 2128 50608 77296
rect 65648 2128 65968 77296
<< obsm4 >>
rect 2083 3027 4128 76941
rect 4608 3027 19488 76941
rect 19968 3027 34848 76941
rect 35328 3027 50208 76941
rect 50688 3027 65568 76941
rect 66048 3027 76666 76941
<< labels >>
rlabel metal2 s 570 0 626 800 6 active
port 1 nsew signal input
rlabel metal3 s 77650 67736 78450 67856 6 io_in[0]
port 2 nsew signal input
rlabel metal2 s 13450 78800 13506 79600 6 io_in[10]
port 3 nsew signal input
rlabel metal2 s 10966 78800 11022 79600 6 io_in[11]
port 4 nsew signal input
rlabel metal2 s 8482 78800 8538 79600 6 io_in[12]
port 5 nsew signal input
rlabel metal2 s 6090 78800 6146 79600 6 io_in[13]
port 6 nsew signal input
rlabel metal3 s 77650 56448 78450 56568 6 io_in[14]
port 7 nsew signal input
rlabel metal3 s 77650 55360 78450 55480 6 io_in[15]
port 8 nsew signal input
rlabel metal2 s 3606 78800 3662 79600 6 io_in[16]
port 9 nsew signal input
rlabel metal2 s 1214 78800 1270 79600 6 io_in[17]
port 10 nsew signal input
rlabel metal3 s 77650 11704 78450 11824 6 io_in[18]
port 11 nsew signal input
rlabel metal3 s 77650 10616 78450 10736 6 io_in[19]
port 12 nsew signal input
rlabel metal3 s 77650 66648 78450 66768 6 io_in[1]
port 13 nsew signal input
rlabel metal3 s 77650 54272 78450 54392 6 io_in[20]
port 14 nsew signal input
rlabel metal3 s 77650 53184 78450 53304 6 io_in[21]
port 15 nsew signal input
rlabel metal3 s 77650 9392 78450 9512 6 io_in[22]
port 16 nsew signal input
rlabel metal3 s 77650 8304 78450 8424 6 io_in[23]
port 17 nsew signal input
rlabel metal3 s 77650 7216 78450 7336 6 io_in[24]
port 18 nsew signal input
rlabel metal3 s 77650 6128 78450 6248 6 io_in[25]
port 19 nsew signal input
rlabel metal3 s 77650 4904 78450 5024 6 io_in[26]
port 20 nsew signal input
rlabel metal3 s 77650 52096 78450 52216 6 io_in[27]
port 21 nsew signal input
rlabel metal3 s 77650 50872 78450 50992 6 io_in[28]
port 22 nsew signal input
rlabel metal3 s 77650 49784 78450 49904 6 io_in[29]
port 23 nsew signal input
rlabel metal3 s 77650 65424 78450 65544 6 io_in[2]
port 24 nsew signal input
rlabel metal3 s 77650 3816 78450 3936 6 io_in[30]
port 25 nsew signal input
rlabel metal3 s 77650 2728 78450 2848 6 io_in[31]
port 26 nsew signal input
rlabel metal3 s 77650 1640 78450 1760 6 io_in[32]
port 27 nsew signal input
rlabel metal3 s 77650 552 78450 672 6 io_in[33]
port 28 nsew signal input
rlabel metal3 s 77650 48696 78450 48816 6 io_in[34]
port 29 nsew signal input
rlabel metal3 s 77650 47608 78450 47728 6 io_in[35]
port 30 nsew signal input
rlabel metal3 s 77650 46384 78450 46504 6 io_in[36]
port 31 nsew signal input
rlabel metal3 s 77650 45296 78450 45416 6 io_in[37]
port 32 nsew signal input
rlabel metal3 s 77650 64336 78450 64456 6 io_in[3]
port 33 nsew signal input
rlabel metal3 s 77650 63248 78450 63368 6 io_in[4]
port 34 nsew signal input
rlabel metal3 s 77650 62160 78450 62280 6 io_in[5]
port 35 nsew signal input
rlabel metal3 s 77650 60936 78450 61056 6 io_in[6]
port 36 nsew signal input
rlabel metal3 s 77650 59848 78450 59968 6 io_in[7]
port 37 nsew signal input
rlabel metal3 s 77650 58760 78450 58880 6 io_in[8]
port 38 nsew signal input
rlabel metal3 s 77650 57672 78450 57792 6 io_in[9]
port 39 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 io_oeb[0]
port 40 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 io_oeb[10]
port 41 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 io_oeb[11]
port 42 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 io_oeb[12]
port 43 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 io_oeb[13]
port 44 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 io_oeb[14]
port 45 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 io_oeb[15]
port 46 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 io_oeb[16]
port 47 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 io_oeb[17]
port 48 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 io_oeb[18]
port 49 nsew signal output
rlabel metal3 s 0 2456 800 2576 6 io_oeb[19]
port 50 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 io_oeb[1]
port 51 nsew signal output
rlabel metal3 s 0 824 800 944 6 io_oeb[20]
port 52 nsew signal output
rlabel metal2 s 77206 78800 77262 79600 6 io_oeb[21]
port 53 nsew signal output
rlabel metal2 s 74722 78800 74778 79600 6 io_oeb[22]
port 54 nsew signal output
rlabel metal2 s 72330 78800 72386 79600 6 io_oeb[23]
port 55 nsew signal output
rlabel metal2 s 69846 78800 69902 79600 6 io_oeb[24]
port 56 nsew signal output
rlabel metal2 s 67362 78800 67418 79600 6 io_oeb[25]
port 57 nsew signal output
rlabel metal2 s 64970 78800 65026 79600 6 io_oeb[26]
port 58 nsew signal output
rlabel metal2 s 62486 78800 62542 79600 6 io_oeb[27]
port 59 nsew signal output
rlabel metal2 s 60002 78800 60058 79600 6 io_oeb[28]
port 60 nsew signal output
rlabel metal2 s 57610 78800 57666 79600 6 io_oeb[29]
port 61 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 io_oeb[2]
port 62 nsew signal output
rlabel metal2 s 55126 78800 55182 79600 6 io_oeb[30]
port 63 nsew signal output
rlabel metal2 s 52642 78800 52698 79600 6 io_oeb[31]
port 64 nsew signal output
rlabel metal2 s 50250 78800 50306 79600 6 io_oeb[32]
port 65 nsew signal output
rlabel metal2 s 47766 78800 47822 79600 6 io_oeb[33]
port 66 nsew signal output
rlabel metal2 s 45282 78800 45338 79600 6 io_oeb[34]
port 67 nsew signal output
rlabel metal2 s 42890 78800 42946 79600 6 io_oeb[35]
port 68 nsew signal output
rlabel metal2 s 40406 78800 40462 79600 6 io_oeb[36]
port 69 nsew signal output
rlabel metal2 s 37922 78800 37978 79600 6 io_oeb[37]
port 70 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 io_oeb[3]
port 71 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 io_oeb[4]
port 72 nsew signal output
rlabel metal3 s 0 26120 800 26240 6 io_oeb[5]
port 73 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 io_oeb[6]
port 74 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 io_oeb[7]
port 75 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 io_oeb[8]
port 76 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 77650 44208 78450 44328 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 77650 32920 78450 33040 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 77650 31832 78450 31952 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 77650 30744 78450 30864 6 io_out[12]
port 81 nsew signal output
rlabel metal3 s 77650 29656 78450 29776 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 77650 28432 78450 28552 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 77650 27344 78450 27464 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 77650 26256 78450 26376 6 io_out[16]
port 85 nsew signal output
rlabel metal3 s 77650 25168 78450 25288 6 io_out[17]
port 86 nsew signal output
rlabel metal3 s 77650 24080 78450 24200 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 77650 22856 78450 22976 6 io_out[19]
port 88 nsew signal output
rlabel metal3 s 77650 43120 78450 43240 6 io_out[1]
port 89 nsew signal output
rlabel metal3 s 77650 21768 78450 21888 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 77650 20680 78450 20800 6 io_out[21]
port 91 nsew signal output
rlabel metal3 s 77650 19592 78450 19712 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 77650 18368 78450 18488 6 io_out[23]
port 93 nsew signal output
rlabel metal3 s 77650 17280 78450 17400 6 io_out[24]
port 94 nsew signal output
rlabel metal3 s 77650 16192 78450 16312 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 77650 15104 78450 15224 6 io_out[26]
port 96 nsew signal output
rlabel metal3 s 77650 13880 78450 14000 6 io_out[27]
port 97 nsew signal output
rlabel metal3 s 77650 12792 78450 12912 6 io_out[28]
port 98 nsew signal output
rlabel metal2 s 35530 78800 35586 79600 6 io_out[29]
port 99 nsew signal output
rlabel metal3 s 77650 41896 78450 42016 6 io_out[2]
port 100 nsew signal output
rlabel metal2 s 33046 78800 33102 79600 6 io_out[30]
port 101 nsew signal output
rlabel metal2 s 30562 78800 30618 79600 6 io_out[31]
port 102 nsew signal output
rlabel metal2 s 28170 78800 28226 79600 6 io_out[32]
port 103 nsew signal output
rlabel metal2 s 25686 78800 25742 79600 6 io_out[33]
port 104 nsew signal output
rlabel metal2 s 23202 78800 23258 79600 6 io_out[34]
port 105 nsew signal output
rlabel metal2 s 20810 78800 20866 79600 6 io_out[35]
port 106 nsew signal output
rlabel metal2 s 18326 78800 18382 79600 6 io_out[36]
port 107 nsew signal output
rlabel metal2 s 15842 78800 15898 79600 6 io_out[37]
port 108 nsew signal output
rlabel metal3 s 77650 40808 78450 40928 6 io_out[3]
port 109 nsew signal output
rlabel metal3 s 77650 39720 78450 39840 6 io_out[4]
port 110 nsew signal output
rlabel metal3 s 77650 38632 78450 38752 6 io_out[5]
port 111 nsew signal output
rlabel metal3 s 77650 37408 78450 37528 6 io_out[6]
port 112 nsew signal output
rlabel metal3 s 77650 36320 78450 36440 6 io_out[7]
port 113 nsew signal output
rlabel metal3 s 77650 35232 78450 35352 6 io_out[8]
port 114 nsew signal output
rlabel metal3 s 77650 34144 78450 34264 6 io_out[9]
port 115 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 la1_data_in[0]
port 116 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la1_data_in[10]
port 117 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la1_data_in[11]
port 118 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 la1_data_in[12]
port 119 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 la1_data_in[13]
port 120 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 la1_data_in[14]
port 121 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 la1_data_in[15]
port 122 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 la1_data_in[16]
port 123 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 la1_data_in[17]
port 124 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 la1_data_in[18]
port 125 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 la1_data_in[19]
port 126 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la1_data_in[1]
port 127 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 la1_data_in[20]
port 128 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 la1_data_in[21]
port 129 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 la1_data_in[22]
port 130 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 la1_data_in[23]
port 131 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 la1_data_in[24]
port 132 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 la1_data_in[25]
port 133 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 la1_data_in[26]
port 134 nsew signal input
rlabel metal3 s 77650 72224 78450 72344 6 la1_data_in[27]
port 135 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 la1_data_in[28]
port 136 nsew signal input
rlabel metal3 s 77650 71136 78450 71256 6 la1_data_in[29]
port 137 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la1_data_in[2]
port 138 nsew signal input
rlabel metal3 s 77650 69912 78450 70032 6 la1_data_in[30]
port 139 nsew signal input
rlabel metal3 s 77650 68824 78450 68944 6 la1_data_in[31]
port 140 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 la1_data_in[3]
port 141 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la1_data_in[4]
port 142 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la1_data_in[5]
port 143 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 la1_data_in[6]
port 144 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la1_data_in[7]
port 145 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 la1_data_in[8]
port 146 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 la1_data_in[9]
port 147 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 la1_data_out[0]
port 148 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la1_data_out[10]
port 149 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la1_data_out[11]
port 150 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la1_data_out[12]
port 151 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la1_data_out[13]
port 152 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la1_data_out[14]
port 153 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 la1_data_out[15]
port 154 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la1_data_out[16]
port 155 nsew signal output
rlabel metal2 s 56230 0 56286 800 6 la1_data_out[17]
port 156 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 la1_data_out[18]
port 157 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la1_data_out[19]
port 158 nsew signal output
rlabel metal2 s 76470 0 76526 800 6 la1_data_out[1]
port 159 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la1_data_out[20]
port 160 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 la1_data_out[21]
port 161 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 la1_data_out[22]
port 162 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 la1_data_out[23]
port 163 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la1_data_out[24]
port 164 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la1_data_out[25]
port 165 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la1_data_out[26]
port 166 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la1_data_out[27]
port 167 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 la1_data_out[28]
port 168 nsew signal output
rlabel metal2 s 41050 0 41106 800 6 la1_data_out[29]
port 169 nsew signal output
rlabel metal2 s 75182 0 75238 800 6 la1_data_out[2]
port 170 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 la1_data_out[30]
port 171 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 la1_data_out[31]
port 172 nsew signal output
rlabel metal2 s 73894 0 73950 800 6 la1_data_out[3]
port 173 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 la1_data_out[4]
port 174 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 la1_data_out[5]
port 175 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 la1_data_out[6]
port 176 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 la1_data_out[7]
port 177 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 la1_data_out[8]
port 178 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 la1_data_out[9]
port 179 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 la1_oenb[0]
port 180 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 la1_oenb[10]
port 181 nsew signal input
rlabel metal3 s 0 59984 800 60104 6 la1_oenb[11]
port 182 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 la1_oenb[12]
port 183 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 la1_oenb[13]
port 184 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 la1_oenb[14]
port 185 nsew signal input
rlabel metal3 s 0 53184 800 53304 6 la1_oenb[15]
port 186 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 la1_oenb[16]
port 187 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 la1_oenb[17]
port 188 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 la1_oenb[18]
port 189 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 la1_oenb[19]
port 190 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 la1_oenb[1]
port 191 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 la1_oenb[20]
port 192 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 la1_oenb[21]
port 193 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 la1_oenb[22]
port 194 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 la1_oenb[23]
port 195 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 la1_oenb[24]
port 196 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 la1_oenb[25]
port 197 nsew signal input
rlabel metal3 s 77650 78888 78450 79008 6 la1_oenb[26]
port 198 nsew signal input
rlabel metal3 s 77650 77800 78450 77920 6 la1_oenb[27]
port 199 nsew signal input
rlabel metal3 s 77650 76712 78450 76832 6 la1_oenb[28]
port 200 nsew signal input
rlabel metal3 s 77650 75624 78450 75744 6 la1_oenb[29]
port 201 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 la1_oenb[2]
port 202 nsew signal input
rlabel metal3 s 77650 74400 78450 74520 6 la1_oenb[30]
port 203 nsew signal input
rlabel metal3 s 77650 73312 78450 73432 6 la1_oenb[31]
port 204 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 la1_oenb[3]
port 205 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 la1_oenb[4]
port 206 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 la1_oenb[5]
port 207 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 la1_oenb[6]
port 208 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 la1_oenb[7]
port 209 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 la1_oenb[8]
port 210 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 la1_oenb[9]
port 211 nsew signal input
rlabel metal4 s 4208 2128 4528 77296 6 vccd1
port 212 nsew power input
rlabel metal4 s 34928 2128 35248 77296 6 vccd1
port 212 nsew power input
rlabel metal4 s 65648 2128 65968 77296 6 vccd1
port 212 nsew power input
rlabel metal4 s 19568 2128 19888 77296 6 vssd1
port 213 nsew ground input
rlabel metal4 s 50288 2128 50608 77296 6 vssd1
port 213 nsew ground input
rlabel metal2 s 1766 0 1822 800 6 wb_clk_i
port 214 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 78450 79600
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 22649010
string GDS_FILE /openlane/designs/wrapped_hack_soc_dffram/runs/RUN_2022.03.16_16.06.18/results/finishing/wrapped_hack_soc_dffram.magic.gds
string GDS_START 14984616
<< end >>

