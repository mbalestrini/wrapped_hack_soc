* NGSPICE file created from wrapped_hack_soc_dffram.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for DFFRF_2R1W abstract view
.subckt DFFRF_2R1W CLK DA[0] DA[10] DA[11] DA[12] DA[13] DA[14] DA[15] DA[16] DA[17]
+ DA[18] DA[19] DA[1] DA[20] DA[21] DA[22] DA[23] DA[24] DA[25] DA[26] DA[27] DA[28]
+ DA[29] DA[2] DA[30] DA[31] DA[3] DA[4] DA[5] DA[6] DA[7] DA[8] DA[9] DB[0] DB[10]
+ DB[11] DB[12] DB[13] DB[14] DB[15] DB[16] DB[17] DB[18] DB[19] DB[1] DB[20] DB[21]
+ DB[22] DB[23] DB[24] DB[25] DB[26] DB[27] DB[28] DB[29] DB[2] DB[30] DB[31] DB[3]
+ DB[4] DB[5] DB[6] DB[7] DB[8] DB[9] DW[0] DW[10] DW[11] DW[12] DW[13] DW[14] DW[15]
+ DW[16] DW[17] DW[18] DW[19] DW[1] DW[20] DW[21] DW[22] DW[23] DW[24] DW[25] DW[26]
+ DW[27] DW[28] DW[29] DW[2] DW[30] DW[31] DW[3] DW[4] DW[5] DW[6] DW[7] DW[8] DW[9]
+ RA[0] RA[1] RA[2] RA[3] RA[4] RB[0] RB[1] RB[2] RB[3] RB[4] RW[0] RW[1] RW[2] RW[3]
+ RW[4] VGND VPWR WE
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt wrapped_hack_soc_dffram active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ vccd1 vssd1 wb_clk_i
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3155_ _3187_/A _3155_/B vssd1 vssd1 vccd1 vccd1 _3155_/X sky130_fd_sc_hd__or2_1
X_3086_ _3154_/A _3086_/B vssd1 vssd1 vccd1 vccd1 _4833_/B sky130_fd_sc_hd__xor2_4
XFILLER_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ _5107_/Q _3983_/X _3980_/A _3186_/X vssd1 vssd1 vccd1 vccd1 _5107_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2939_ _2939_/A _2939_/B vssd1 vssd1 vccd1 vccd1 _2939_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_2_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4609_ _4609_/A _4609_/B vssd1 vssd1 vccd1 vccd1 _4610_/A sky130_fd_sc_hd__and2_1
X_5589_ _5589_/A _2619_/Y vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__ebufn_8
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4960_ _4958_/Y _4959_/X _2787_/B vssd1 vssd1 vccd1 vccd1 _5445_/D sky130_fd_sc_hd__a21oi_1
X_4891_ _5383_/D _4884_/X _4890_/Y _4882_/X vssd1 vssd1 vccd1 vccd1 _5415_/D sky130_fd_sc_hd__o211a_1
X_3911_ _3911_/A vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__clkbuf_2
X_3842_ _3841_/B _3835_/A _3834_/A _3841_/A vssd1 vssd1 vccd1 vccd1 _3843_/C sky130_fd_sc_hd__a31o_1
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3773_ _3773_/A0 _3773_/A1 _3773_/S vssd1 vssd1 vccd1 vccd1 _3773_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2724_ _5037_/Q _5040_/Q vssd1 vssd1 vccd1 vccd1 _2725_/B sky130_fd_sc_hd__or2_1
X_5443_ _5443_/CLK _5443_/D vssd1 vssd1 vccd1 vccd1 _5443_/Q sky130_fd_sc_hd__dfxtp_1
X_2655_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2655_/Y sky130_fd_sc_hd__inv_2
X_5374_ _5403_/Q _5374_/D vssd1 vssd1 vccd1 vccd1 _5374_/Q sky130_fd_sc_hd__dfxtp_1
X_2586_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2591_/A sky130_fd_sc_hd__buf_6
X_4325_ _4325_/A vssd1 vssd1 vccd1 vccd1 _5222_/D sky130_fd_sc_hd__clkbuf_1
X_4256_ _4609_/A _4256_/B vssd1 vssd1 vccd1 vccd1 _4257_/A sky130_fd_sc_hd__and2_1
XFILLER_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3207_ _3275_/A _3207_/B vssd1 vssd1 vccd1 vccd1 _3224_/A sky130_fd_sc_hd__or2_1
X_4187_ _5409_/Q _5360_/Q _4199_/S vssd1 vssd1 vccd1 vccd1 _4187_/X sky130_fd_sc_hd__mux2_1
X_3138_ _3647_/A _5399_/Q vssd1 vssd1 vccd1 vccd1 _3139_/B sky130_fd_sc_hd__and2_1
XFILLER_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3069_ _3126_/B vssd1 vssd1 vccd1 vccd1 _3139_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4110_ hold37/A _4109_/A _4094_/X vssd1 vssd1 vccd1 vccd1 _4110_/Y sky130_fd_sc_hd__a21oi_1
X_5090_ _5323_/CLK _5090_/D vssd1 vssd1 vccd1 vccd1 _5090_/Q sky130_fd_sc_hd__dfxtp_1
X_4041_ _3462_/B _4041_/B vssd1 vssd1 vccd1 vccd1 _4042_/B sky130_fd_sc_hd__and2b_1
XFILLER_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4943_ _4943_/A vssd1 vssd1 vccd1 vccd1 _5438_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4874_ _5379_/D _4863_/X _4873_/Y _4861_/X vssd1 vssd1 vccd1 vccd1 _5411_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3825_ _3758_/X _3823_/X _3824_/X _3698_/A vssd1 vssd1 vccd1 vccd1 _3838_/A sky130_fd_sc_hd__o31a_1
XFILLER_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3756_ _3755_/X _5026_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3757_/A sky130_fd_sc_hd__mux2_1
X_2707_ _5117_/Q _5116_/Q _5115_/Q _5114_/Q vssd1 vssd1 vccd1 vccd1 _2752_/B sky130_fd_sc_hd__or4_4
X_5426_ _5430_/CLK _5426_/D vssd1 vssd1 vccd1 vccd1 _5426_/Q sky130_fd_sc_hd__dfxtp_1
X_3687_ _5323_/Q _4587_/B _4328_/B vssd1 vssd1 vccd1 vccd1 _4589_/A sky130_fd_sc_hd__and3_1
X_2638_ _2640_/A vssd1 vssd1 vccd1 vccd1 _2638_/Y sky130_fd_sc_hd__inv_2
X_5357_ _5444_/CLK _5357_/D vssd1 vssd1 vccd1 vccd1 _5357_/Q sky130_fd_sc_hd__dfxtp_1
X_2569_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2569_/Y sky130_fd_sc_hd__inv_2
X_4308_ _5214_/Q _4264_/X _4307_/X vssd1 vssd1 vccd1 vccd1 _4308_/X sky130_fd_sc_hd__a21o_1
X_5288_ _5435_/CLK _5288_/D vssd1 vssd1 vccd1 vccd1 _5288_/Q sky130_fd_sc_hd__dfxtp_1
X_4239_ _5200_/Q _5196_/Q _4251_/S vssd1 vssd1 vccd1 vccd1 _4240_/B sky130_fd_sc_hd__mux2_1
XFILLER_28_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3610_ _4504_/A vssd1 vssd1 vccd1 vccd1 _4594_/A sky130_fd_sc_hd__clkbuf_2
X_4590_ _4589_/Y _4330_/X _4692_/C vssd1 vssd1 vccd1 vccd1 _4591_/B sky130_fd_sc_hd__a21o_1
X_3541_ _4285_/A vssd1 vssd1 vccd1 vccd1 _3541_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_6_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3472_ _3472_/A _3472_/B vssd1 vssd1 vccd1 vccd1 _4038_/B sky130_fd_sc_hd__and2_1
X_5211_ _5369_/CLK _5211_/D vssd1 vssd1 vccd1 vccd1 _5211_/Q sky130_fd_sc_hd__dfxtp_1
X_5142_ _5313_/CLK _5142_/D vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
X_5073_ _5077_/CLK _5073_/D vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfxtp_1
X_4024_ _4024_/A _4024_/B vssd1 vssd1 vccd1 vccd1 _4033_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4926_ _4926_/A vssd1 vssd1 vccd1 vccd1 _5428_/D sky130_fd_sc_hd__clkbuf_1
X_4857_ _5375_/D _4840_/X _4856_/Y _4842_/X vssd1 vssd1 vccd1 vccd1 _5407_/D sky130_fd_sc_hd__o211a_1
X_3808_ _5047_/Q _3810_/C _3800_/X vssd1 vssd1 vccd1 vccd1 _3809_/B sky130_fd_sc_hd__o21ai_1
XFILLER_20_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4788_ _5336_/Q _4945_/C _5370_/Q vssd1 vssd1 vccd1 vccd1 _4789_/C sky130_fd_sc_hd__mux2_1
X_3739_ _3739_/A vssd1 vssd1 vccd1 vccd1 _5023_/D sky130_fd_sc_hd__clkbuf_1
X_5409_ _5403_/Q _5409_/D vssd1 vssd1 vccd1 vccd1 _5409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5521__111 vssd1 vssd1 vccd1 vccd1 _5521__111/HI _5637_/A sky130_fd_sc_hd__conb_1
XFILLER_0_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2972_ _3033_/A vssd1 vssd1 vccd1 vccd1 _3130_/A sky130_fd_sc_hd__buf_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4711_ _4711_/A vssd1 vssd1 vccd1 vccd1 _5329_/D sky130_fd_sc_hd__clkbuf_1
X_4642_ _4642_/A vssd1 vssd1 vccd1 vccd1 _5312_/D sky130_fd_sc_hd__clkbuf_1
X_4573_ _5296_/Q _4577_/B vssd1 vssd1 vccd1 vccd1 _4573_/X sky130_fd_sc_hd__or2_1
X_3524_ _3524_/A vssd1 vssd1 vccd1 vccd1 _3682_/C sky130_fd_sc_hd__clkbuf_1
X_3455_ _4022_/A _4042_/A _3455_/C vssd1 vssd1 vccd1 vccd1 _3455_/X sky130_fd_sc_hd__or3_1
X_3386_ _3338_/A _3382_/X _3385_/Y _3344_/X vssd1 vssd1 vccd1 vccd1 _3387_/C sky130_fd_sc_hd__a211o_1
X_5125_ _5126_/CLK _5125_/D vssd1 vssd1 vccd1 vccd1 _5125_/Q sky130_fd_sc_hd__dfxtp_1
X_5056_ _5058_/CLK _5056_/D vssd1 vssd1 vccd1 vccd1 _5056_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4909_ _5420_/Q _4908_/Y _5437_/D vssd1 vssd1 vccd1 vccd1 _5420_/D sky130_fd_sc_hd__a21o_1
XFILLER_5_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_14_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5437_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_5 _5640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3252_/S _3240_/B vssd1 vssd1 vccd1 vccd1 _3240_/Y sky130_fd_sc_hd__nand2_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3187_/A _5241_/Q vssd1 vssd1 vccd1 vccd1 _3171_/X sky130_fd_sc_hd__or2_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2955_ input40/X _2952_/Y _2953_/X _2954_/X vssd1 vssd1 vccd1 vccd1 _2955_/X sky130_fd_sc_hd__a211o_1
XFILLER_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2886_ _5238_/Q _2886_/B vssd1 vssd1 vccd1 vccd1 _2913_/A sky130_fd_sc_hd__xnor2_1
X_4625_ _4625_/A vssd1 vssd1 vccd1 vccd1 _5308_/D sky130_fd_sc_hd__clkbuf_1
X_4556_ input2/X _4552_/X _4555_/X _4416_/X vssd1 vssd1 vccd1 vccd1 _5289_/D sky130_fd_sc_hd__o211a_1
X_3507_ _5251_/Q vssd1 vssd1 vccd1 vccd1 _3510_/A sky130_fd_sc_hd__inv_2
X_4487_ _4487_/A vssd1 vssd1 vccd1 vccd1 _5263_/D sky130_fd_sc_hd__clkbuf_1
X_3438_ _3572_/A _3438_/B vssd1 vssd1 vccd1 vccd1 _3439_/D sky130_fd_sc_hd__nor2_1
X_3369_ _3393_/A _3353_/X _3393_/B _3368_/X vssd1 vssd1 vccd1 vccd1 _3369_/Y sky130_fd_sc_hd__a211oi_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _5436_/CLK _5108_/D vssd1 vssd1 vccd1 vccd1 _5108_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5039_ _5439_/CLK _5039_/D vssd1 vssd1 vccd1 vccd1 _5039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2740_ _5037_/Q vssd1 vssd1 vccd1 vccd1 _3754_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2671_ _2671_/A vssd1 vssd1 vccd1 vccd1 _2671_/Y sky130_fd_sc_hd__inv_2
X_4410_ _5239_/Q _4402_/X _4409_/X _4397_/X vssd1 vssd1 vccd1 vccd1 _5239_/D sky130_fd_sc_hd__o211a_1
X_5390_ _5403_/Q _5390_/D vssd1 vssd1 vccd1 vccd1 _5390_/Q sky130_fd_sc_hd__dfxtp_1
X_4341_ _4341_/A vssd1 vssd1 vccd1 vccd1 _5224_/D sky130_fd_sc_hd__clkbuf_1
X_4272_ _5186_/Q _3682_/D _4275_/A _5008_/Q vssd1 vssd1 vccd1 vccd1 _4272_/X sky130_fd_sc_hd__a22o_1
X_3223_ _3223_/A _3223_/B vssd1 vssd1 vccd1 vccd1 _3240_/B sky130_fd_sc_hd__nor2_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3154_ _3154_/A _3154_/B vssd1 vssd1 vccd1 vccd1 _4834_/C sky130_fd_sc_hd__xnor2_4
X_3085_ _3118_/S _3081_/Y _3102_/B _3084_/Y vssd1 vssd1 vccd1 vccd1 _3086_/B sky130_fd_sc_hd__a31o_1
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3987_ _5106_/Q _3983_/X _3980_/A _3170_/X vssd1 vssd1 vccd1 vccd1 _5106_/D sky130_fd_sc_hd__a22o_1
X_2938_ _2938_/A _2938_/B vssd1 vssd1 vccd1 vccd1 _2939_/B sky130_fd_sc_hd__nand2_1
XFILLER_136_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2869_ _2869_/A _4999_/Q vssd1 vssd1 vccd1 vccd1 _2869_/X sky130_fd_sc_hd__and2_1
X_4608_ _5305_/Q _4607_/X _4617_/S vssd1 vssd1 vccd1 vccd1 _4609_/B sky130_fd_sc_hd__mux2_1
X_5588_ _5588_/A _2618_/Y vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__ebufn_8
X_4539_ _5283_/Q _5430_/Q _4541_/S vssd1 vssd1 vccd1 vccd1 _4540_/A sky130_fd_sc_hd__mux2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4890_ _4893_/B _4889_/Y _4841_/B vssd1 vssd1 vccd1 vccd1 _4890_/Y sky130_fd_sc_hd__o21ai_1
X_3910_ _3910_/A vssd1 vssd1 vccd1 vccd1 _3910_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3841_ _3841_/A _3841_/B _3847_/C vssd1 vssd1 vccd1 vccd1 _3841_/X sky130_fd_sc_hd__and3_1
X_3772_ _3823_/B _3772_/B vssd1 vssd1 vccd1 vccd1 _3772_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2723_ _5039_/Q vssd1 vssd1 vccd1 vccd1 _2753_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5442_ _5443_/CLK _5442_/D vssd1 vssd1 vccd1 vccd1 _5442_/Q sky130_fd_sc_hd__dfxtp_1
X_2654_ _2666_/A vssd1 vssd1 vccd1 vccd1 _2659_/A sky130_fd_sc_hd__buf_2
X_5373_ _5403_/Q _5373_/D vssd1 vssd1 vccd1 vccd1 _5373_/Q sky130_fd_sc_hd__dfxtp_1
X_2585_ _2585_/A vssd1 vssd1 vccd1 vccd1 _2585_/Y sky130_fd_sc_hd__inv_2
X_4324_ _4323_/X _5222_/Q _4324_/S vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4255_ _5205_/Q _5201_/Q _4258_/S vssd1 vssd1 vccd1 vccd1 _4256_/B sky130_fd_sc_hd__mux2_1
X_3206_ _3402_/A _3829_/A _3823_/D _3284_/A _3205_/Y vssd1 vssd1 vccd1 vccd1 _3207_/B
+ sky130_fd_sc_hd__a41o_1
X_4186_ _4203_/A vssd1 vssd1 vccd1 vccd1 _4199_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3137_ _5383_/Q _3028_/A _4833_/C _3120_/X _3136_/X vssd1 vssd1 vccd1 vccd1 _5383_/D
+ sky130_fd_sc_hd__o221a_1
X_3068_ _3036_/A _3056_/X _3067_/C _3038_/X _3066_/C vssd1 vssd1 vccd1 vccd1 _3081_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5500__90 vssd1 vssd1 vccd1 vccd1 _5500__90/HI _5599_/A sky130_fd_sc_hd__conb_1
XFILLER_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4040_ _2838_/X _4030_/Y _4039_/X _4025_/Y vssd1 vssd1 vccd1 vccd1 _5131_/D sky130_fd_sc_hd__a211o_1
XFILLER_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4942_ _4829_/S _5227_/Q _5419_/Q _4942_/D vssd1 vssd1 vccd1 vccd1 _4943_/A sky130_fd_sc_hd__and4b_1
X_4873_ _4901_/A _4873_/B vssd1 vssd1 vccd1 vccd1 _4873_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3824_ _3851_/A _3824_/B _3824_/C _3853_/A vssd1 vssd1 vccd1 vccd1 _3824_/X sky130_fd_sc_hd__or4b_1
X_3755_ _3749_/Y _3750_/X _3751_/Y _3753_/X _3754_/X vssd1 vssd1 vccd1 vccd1 _3755_/X
+ sky130_fd_sc_hd__a32o_1
X_3686_ _5010_/Q _4266_/S _3682_/X _5180_/Q vssd1 vssd1 vccd1 vccd1 _5010_/D sky130_fd_sc_hd__a22o_1
X_2706_ _2706_/A _2706_/B vssd1 vssd1 vccd1 vccd1 _2706_/Y sky130_fd_sc_hd__nor2_1
X_2637_ _2640_/A vssd1 vssd1 vccd1 vccd1 _2637_/Y sky130_fd_sc_hd__inv_2
X_5425_ _5430_/CLK _5425_/D vssd1 vssd1 vccd1 vccd1 _5425_/Q sky130_fd_sc_hd__dfxtp_1
X_5356_ _5444_/CLK _5356_/D vssd1 vssd1 vccd1 vccd1 _5356_/Q sky130_fd_sc_hd__dfxtp_1
X_2568_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2568_/Y sky130_fd_sc_hd__inv_2
X_4307_ _5168_/Q _4285_/A _4276_/A _5194_/Q vssd1 vssd1 vccd1 vccd1 _4307_/X sky130_fd_sc_hd__a22o_1
X_5287_ _5435_/CLK _5287_/D vssd1 vssd1 vccd1 vccd1 _5287_/Q sky130_fd_sc_hd__dfxtp_1
X_4238_ _4258_/S vssd1 vssd1 vccd1 vccd1 _4251_/S sky130_fd_sc_hd__clkbuf_2
X_4169_ _4203_/A vssd1 vssd1 vccd1 vccd1 _4182_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5477__67 vssd1 vssd1 vccd1 vccd1 _5477__67/HI _5554_/A sky130_fd_sc_hd__conb_1
XFILLER_46_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3540_ _5583_/A _3677_/B _3539_/X _2761_/X vssd1 vssd1 vccd1 vccd1 _4984_/D sky130_fd_sc_hd__a211o_1
XFILLER_10_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5210_ _5339_/CLK _5210_/D vssd1 vssd1 vccd1 vccd1 _5210_/Q sky130_fd_sc_hd__dfxtp_1
X_3471_ _3464_/B _2822_/B _2838_/A vssd1 vssd1 vccd1 vccd1 _3472_/B sky130_fd_sc_hd__o21ai_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5141_ _5313_/CLK _5141_/D vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dfxtp_1
X_5072_ _5077_/CLK _5072_/D vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
X_4023_ _3773_/S _2725_/B _2744_/B _3754_/A _3726_/B vssd1 vssd1 vccd1 vccd1 _4024_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5491__81 vssd1 vssd1 vccd1 vccd1 _5491__81/HI _5569_/A sky130_fd_sc_hd__conb_1
XFILLER_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4925_ _5428_/Q _5379_/Q _4927_/S vssd1 vssd1 vccd1 vccd1 _4926_/A sky130_fd_sc_hd__mux2_1
X_4856_ _4864_/C _4855_/Y _4851_/X vssd1 vssd1 vccd1 vccd1 _4856_/Y sky130_fd_sc_hd__o21ai_1
X_3807_ _5047_/Q _3810_/C vssd1 vssd1 vccd1 vccd1 _3809_/A sky130_fd_sc_hd__and2_1
X_4787_ hold137/X _4785_/A _4786_/Y vssd1 vssd1 vccd1 vccd1 _5369_/D sky130_fd_sc_hd__a21oi_1
X_3738_ _3737_/X _5023_/Q _3767_/A vssd1 vssd1 vccd1 vccd1 _3739_/A sky130_fd_sc_hd__mux2_1
X_3669_ _5005_/Q _5006_/Q vssd1 vssd1 vccd1 vccd1 _3669_/Y sky130_fd_sc_hd__xnor2_1
X_5408_ _5403_/Q _5408_/D vssd1 vssd1 vccd1 vccd1 _5408_/Q sky130_fd_sc_hd__dfxtp_1
X_5339_ _5339_/CLK _5339_/D vssd1 vssd1 vccd1 vccd1 _5339_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2971_ _3051_/A _2971_/B vssd1 vssd1 vccd1 vccd1 _2984_/A sky130_fd_sc_hd__xnor2_1
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4710_ _4714_/A _4710_/B vssd1 vssd1 vccd1 vccd1 _4711_/A sky130_fd_sc_hd__and2b_1
XFILLER_42_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4641_ _4655_/A _4641_/B vssd1 vssd1 vccd1 vccd1 _4642_/A sky130_fd_sc_hd__and2_1
X_4572_ _5291_/Q _4566_/X _4570_/X _4571_/X vssd1 vssd1 vccd1 vccd1 _5295_/D sky130_fd_sc_hd__o211a_1
X_3523_ _3592_/A vssd1 vssd1 vccd1 vccd1 _3682_/B sky130_fd_sc_hd__clkbuf_1
X_3454_ _3480_/B _3452_/X _3453_/X vssd1 vssd1 vccd1 vccd1 _3455_/C sky130_fd_sc_hd__a21oi_1
X_3385_ _3378_/B _3384_/X _3393_/A vssd1 vssd1 vccd1 vccd1 _3385_/Y sky130_fd_sc_hd__o21ai_1
X_5124_ _5126_/CLK _5124_/D vssd1 vssd1 vccd1 vccd1 _5124_/Q sky130_fd_sc_hd__dfxtp_1
X_5055_ _5439_/CLK _5055_/D vssd1 vssd1 vccd1 vccd1 _5055_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4908_ _4916_/S vssd1 vssd1 vccd1 vccd1 _4908_/Y sky130_fd_sc_hd__inv_2
X_4839_ _4844_/A vssd1 vssd1 vccd1 vccd1 _4841_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__clkbuf_2
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5528__118 vssd1 vssd1 vccd1 vccd1 _5528__118/HI _5528__118/LO sky130_fd_sc_hd__conb_1
XANTENNA_6 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _4835_/A vssd1 vssd1 vccd1 vccd1 _3170_/X sky130_fd_sc_hd__buf_2
XFILLER_47_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5461__51 vssd1 vssd1 vccd1 vccd1 _5461__51/HI _5538_/A sky130_fd_sc_hd__conb_1
XFILLER_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2954_ _5305_/Q _2890_/A _4964_/A _5602_/A _2892_/A vssd1 vssd1 vccd1 vccd1 _2954_/X
+ sky130_fd_sc_hd__a221o_1
X_2885_ _3029_/A _5387_/Q vssd1 vssd1 vccd1 vccd1 _2886_/B sky130_fd_sc_hd__nand2_1
X_4624_ _4632_/A _4624_/B vssd1 vssd1 vccd1 vccd1 _4625_/A sky130_fd_sc_hd__and2_1
X_4555_ _5289_/Q _4564_/B vssd1 vssd1 vccd1 vccd1 _4555_/X sky130_fd_sc_hd__or2_1
X_3506_ _5248_/Q vssd1 vssd1 vccd1 vccd1 _4434_/A sky130_fd_sc_hd__clkbuf_2
X_4486_ _5263_/Q _5101_/Q _4492_/S vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__mux2_1
X_3437_ _3572_/A _3572_/B _3551_/C vssd1 vssd1 vccd1 vccd1 _3578_/B sky130_fd_sc_hd__and3_1
X_3368_ _3352_/S _3366_/Y _3367_/Y _3340_/Y vssd1 vssd1 vccd1 vccd1 _3368_/X sky130_fd_sc_hd__o211a_1
XFILLER_58_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _5437_/CLK _5107_/D vssd1 vssd1 vccd1 vccd1 _5107_/Q sky130_fd_sc_hd__dfxtp_1
X_3299_ _3411_/A _3411_/B vssd1 vssd1 vccd1 vccd1 _3319_/A sky130_fd_sc_hd__or2_1
XFILLER_26_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5038_ _5439_/CLK _5038_/D vssd1 vssd1 vccd1 vccd1 _5038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2670_ _2671_/A vssd1 vssd1 vccd1 vccd1 _2670_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4340_ _4348_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4341_/A sky130_fd_sc_hd__or2_1
X_4271_ _4271_/A vssd1 vssd1 vccd1 vccd1 _5209_/D sky130_fd_sc_hd__clkbuf_1
X_3222_ _3221_/A _3221_/C _3221_/B vssd1 vssd1 vccd1 vccd1 _3223_/B sky130_fd_sc_hd__a21oi_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3153_ _3118_/S _3166_/A _3152_/X vssd1 vssd1 vccd1 vccd1 _3154_/B sky130_fd_sc_hd__o21a_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3084_ _3084_/A _3115_/A vssd1 vssd1 vccd1 vccd1 _3084_/Y sky130_fd_sc_hd__nor2_1
XFILLER_35_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3986_ _5105_/Q _3983_/X _3980_/X _4834_/C vssd1 vssd1 vccd1 vccd1 _5105_/D sky130_fd_sc_hd__a22o_1
X_4004__11 _4005__12/A vssd1 vssd1 vccd1 vccd1 _5118_/CLK sky130_fd_sc_hd__inv_2
X_2937_ _2948_/B _2948_/C _2948_/A vssd1 vssd1 vccd1 vccd1 _2938_/B sky130_fd_sc_hd__a21o_1
X_2868_ _5032_/Q _5031_/Q _2872_/S vssd1 vssd1 vccd1 vccd1 _2868_/X sky130_fd_sc_hd__mux2_1
X_4607_ input4/X _5257_/Q _4616_/S vssd1 vssd1 vccd1 vccd1 _4607_/X sky130_fd_sc_hd__mux2_1
X_2799_ _2870_/A _2870_/B vssd1 vssd1 vccd1 vccd1 _3476_/A sky130_fd_sc_hd__and2_2
X_5587_ _5587_/A _2616_/Y vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__ebufn_8
X_4538_ _4538_/A vssd1 vssd1 vccd1 vccd1 _5282_/D sky130_fd_sc_hd__clkbuf_1
X_4469_ _5256_/Q _5094_/Q _4583_/B vssd1 vssd1 vccd1 vccd1 _4470_/A sky130_fd_sc_hd__mux2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ _3841_/B _3847_/C _3839_/Y vssd1 vssd1 vccd1 vccd1 _5056_/D sky130_fd_sc_hd__o21a_1
XFILLER_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3771_ _5029_/Q _3767_/X _3740_/X _3770_/X vssd1 vssd1 vccd1 vccd1 _5029_/D sky130_fd_sc_hd__a22o_1
X_2722_ _5149_/Q _2727_/A vssd1 vssd1 vccd1 vccd1 _2760_/C sky130_fd_sc_hd__and2_1
XFILLER_8_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5441_ _5443_/CLK _5441_/D vssd1 vssd1 vccd1 vccd1 _5441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2653_ _2653_/A vssd1 vssd1 vccd1 vccd1 _2653_/Y sky130_fd_sc_hd__inv_2
X_2584_ _2585_/A vssd1 vssd1 vccd1 vccd1 _2584_/Y sky130_fd_sc_hd__inv_2
X_5372_ _5403_/Q _5372_/D vssd1 vssd1 vccd1 vccd1 _5372_/Q sky130_fd_sc_hd__dfxtp_1
X_4323_ _5218_/Q _3535_/X _3537_/X _5172_/Q _3543_/B vssd1 vssd1 vccd1 vccd1 _4323_/X
+ sky130_fd_sc_hd__a221o_1
X_4254_ _4611_/A vssd1 vssd1 vccd1 vccd1 _4609_/A sky130_fd_sc_hd__clkbuf_2
X_3205_ _5056_/Q _5057_/Q _3424_/A _5059_/Q vssd1 vssd1 vccd1 vccd1 _3205_/Y sky130_fd_sc_hd__nand4b_1
X_4185_ _4185_/A vssd1 vssd1 vccd1 vccd1 _5184_/D sky130_fd_sc_hd__clkbuf_1
X_3136_ _3187_/A _5239_/Q vssd1 vssd1 vccd1 vccd1 _3136_/X sky130_fd_sc_hd__or2_1
X_3067_ _3067_/A _3067_/B _3067_/C _3005_/A vssd1 vssd1 vccd1 vccd1 _3081_/A sky130_fd_sc_hd__or4b_2
XFILLER_42_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3969_ _5093_/Q _3966_/X _5437_/D _2918_/X vssd1 vssd1 vccd1 vccd1 _5093_/D sky130_fd_sc_hd__a22o_1
X_5639_ _5639_/A _2679_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[35] sky130_fd_sc_hd__ebufn_8
XFILLER_136_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4941_ _4941_/A vssd1 vssd1 vccd1 vccd1 _5435_/D sky130_fd_sc_hd__clkbuf_1
X_4872_ _5411_/Q _4875_/C vssd1 vssd1 vccd1 vccd1 _4873_/B sky130_fd_sc_hd__xnor2_1
Xclkbuf_1_1_0__1653_ clkbuf_0__1653_/X vssd1 vssd1 vccd1 vccd1 _4005__12/A sky130_fd_sc_hd__clkbuf_2
X_3823_ _3823_/A _3823_/B _3829_/A _3823_/D vssd1 vssd1 vccd1 vccd1 _3823_/X sky130_fd_sc_hd__or4_1
XFILLER_32_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_9_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5077_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3754_ _3754_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _3754_/X sky130_fd_sc_hd__and2_1
X_3685_ _5009_/Q _4266_/S _3682_/X _5181_/Q vssd1 vssd1 vccd1 vccd1 _5009_/D sky130_fd_sc_hd__a22o_1
X_2705_ _5050_/Q _5049_/Q _5051_/Q _2705_/D vssd1 vssd1 vccd1 vccd1 _2706_/B sky130_fd_sc_hd__or4_2
X_2636_ _2640_/A vssd1 vssd1 vccd1 vccd1 _2636_/Y sky130_fd_sc_hd__inv_2
X_5424_ _5430_/CLK _5424_/D vssd1 vssd1 vccd1 vccd1 _5424_/Q sky130_fd_sc_hd__dfxtp_1
X_5355_ _5444_/CLK _5355_/D vssd1 vssd1 vccd1 vccd1 _5355_/Q sky130_fd_sc_hd__dfxtp_1
X_2567_ _2698_/A vssd1 vssd1 vccd1 vccd1 _2572_/A sky130_fd_sc_hd__clkbuf_2
X_4306_ _4306_/A vssd1 vssd1 vccd1 vccd1 _5217_/D sky130_fd_sc_hd__clkbuf_1
X_5286_ _5435_/CLK _5286_/D vssd1 vssd1 vccd1 vccd1 _5286_/Q sky130_fd_sc_hd__dfxtp_1
X_4237_ _4611_/A vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4168_ _5179_/Q _4164_/A _4167_/Y vssd1 vssd1 vccd1 vccd1 _5179_/D sky130_fd_sc_hd__a21o_1
X_4099_ hold88/A _4101_/C _4081_/X vssd1 vssd1 vccd1 vccd1 _4100_/B sky130_fd_sc_hd__o21ai_1
X_3119_ _3154_/A _3119_/B vssd1 vssd1 vccd1 vccd1 _4834_/B sky130_fd_sc_hd__xnor2_4
XFILLER_24_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3470_ _4034_/B _3470_/B vssd1 vssd1 vccd1 vccd1 _3470_/Y sky130_fd_sc_hd__xnor2_1
X_5140_ _5313_/CLK _5140_/D vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5071_ _5077_/CLK _5071_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
X_4022_ _4022_/A _4022_/B vssd1 vssd1 vccd1 vccd1 _4022_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4924_ _4924_/A vssd1 vssd1 vccd1 vccd1 _5427_/D sky130_fd_sc_hd__clkbuf_1
X_4855_ _5407_/Q _4855_/B vssd1 vssd1 vccd1 vccd1 _4855_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4786_ _5369_/Q _4785_/A _4742_/X vssd1 vssd1 vccd1 vccd1 _4786_/Y sky130_fd_sc_hd__o21ai_1
X_3806_ _3806_/A vssd1 vssd1 vccd1 vccd1 _5046_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3737_ _3737_/A1 _3734_/B _3754_/B _3736_/Y vssd1 vssd1 vccd1 vccd1 _3737_/X sky130_fd_sc_hd__a31o_1
X_3668_ _4276_/A vssd1 vssd1 vccd1 vccd1 _3682_/D sky130_fd_sc_hd__buf_2
X_5407_ _5403_/Q _5407_/D vssd1 vssd1 vccd1 vccd1 _5407_/Q sky130_fd_sc_hd__dfxtp_1
X_2619_ _2622_/A vssd1 vssd1 vccd1 vccd1 _2619_/Y sky130_fd_sc_hd__inv_2
X_3599_ _2753_/A _3596_/A _3597_/X _3750_/B vssd1 vssd1 vccd1 vccd1 _3733_/B sky130_fd_sc_hd__o31ai_2
X_5338_ _5339_/CLK _5338_/D vssd1 vssd1 vccd1 vccd1 _5338_/Q sky130_fd_sc_hd__dfxtp_1
X_5269_ _5437_/CLK _5269_/D vssd1 vssd1 vccd1 vccd1 _5269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2970_ _3108_/A _5390_/Q vssd1 vssd1 vccd1 vccd1 _2971_/B sky130_fd_sc_hd__and2_1
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4640_ _5312_/Q _4639_/X _4640_/S vssd1 vssd1 vccd1 vccd1 _4641_/B sky130_fd_sc_hd__mux2_1
XFILLER_30_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4571_ _4571_/A vssd1 vssd1 vccd1 vccd1 _4571_/X sky130_fd_sc_hd__clkbuf_2
X_3522_ _3592_/A _3524_/A vssd1 vssd1 vccd1 vccd1 _3677_/B sky130_fd_sc_hd__nand2_1
X_3453_ _2864_/X _2873_/X _2872_/X _2866_/X _3448_/Y vssd1 vssd1 vccd1 vccd1 _3453_/X
+ sky130_fd_sc_hd__a221o_1
X_3384_ _3551_/B _3357_/X _3383_/X _3338_/A vssd1 vssd1 vccd1 vccd1 _3384_/X sky130_fd_sc_hd__o22a_1
X_5123_ _5126_/CLK _5123_/D vssd1 vssd1 vccd1 vccd1 _5123_/Q sky130_fd_sc_hd__dfxtp_1
X_5054_ _5439_/CLK _5054_/D vssd1 vssd1 vccd1 vccd1 _5054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4907_ _4940_/S vssd1 vssd1 vccd1 vccd1 _4916_/S sky130_fd_sc_hd__clkbuf_2
X_4838_ _3656_/Y _4835_/X _4836_/Y _4837_/X _2924_/A vssd1 vssd1 vccd1 vccd1 _4844_/A
+ sky130_fd_sc_hd__a311o_1
X_4769_ _5363_/Q _4771_/C _4762_/X vssd1 vssd1 vccd1 vccd1 _4770_/B sky130_fd_sc_hd__o21ai_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_7 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_23_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5445_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2953_ _5453_/Q _2953_/B _2953_/C vssd1 vssd1 vccd1 vccd1 _2953_/X sky130_fd_sc_hd__and3_1
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5511__101 vssd1 vssd1 vccd1 vccd1 _5511__101/HI _5618_/A sky130_fd_sc_hd__conb_1
X_2884_ _2950_/A vssd1 vssd1 vccd1 vccd1 _3029_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4623_ _5308_/Q _4621_/X _4640_/S vssd1 vssd1 vccd1 vccd1 _4624_/B sky130_fd_sc_hd__mux2_1
X_4554_ _4581_/B vssd1 vssd1 vccd1 vccd1 _4564_/B sky130_fd_sc_hd__clkbuf_1
X_3505_ _4432_/A _3528_/A vssd1 vssd1 vccd1 vccd1 _3592_/A sky130_fd_sc_hd__nand2_1
X_4485_ _4485_/A vssd1 vssd1 vccd1 vccd1 _5262_/D sky130_fd_sc_hd__clkbuf_1
X_3436_ _4073_/B vssd1 vssd1 vccd1 vccd1 _3572_/A sky130_fd_sc_hd__clkbuf_1
X_3367_ _3393_/A vssd1 vssd1 vccd1 vccd1 _3367_/Y sky130_fd_sc_hd__inv_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _5437_/CLK _5106_/D vssd1 vssd1 vccd1 vccd1 _5106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3298_ _3298_/A _3553_/A vssd1 vssd1 vccd1 vccd1 _3411_/B sky130_fd_sc_hd__xnor2_1
X_5037_ _5439_/CLK _5037_/D vssd1 vssd1 vccd1 vccd1 _5037_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5507__97 vssd1 vssd1 vccd1 vccd1 _5507__97/HI _5610_/A sky130_fd_sc_hd__conb_1
XFILLER_1_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4270_ _4268_/X _5209_/Q _4288_/S vssd1 vssd1 vccd1 vccd1 _4271_/A sky130_fd_sc_hd__mux2_1
X_3221_ _3221_/A _3221_/B _3221_/C vssd1 vssd1 vccd1 vccd1 _3223_/A sky130_fd_sc_hd__and3_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3152_ _3152_/A _3646_/A _3166_/B vssd1 vssd1 vccd1 vccd1 _3152_/X sky130_fd_sc_hd__or3b_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3083_ _3083_/A _3083_/B vssd1 vssd1 vccd1 vccd1 _3115_/A sky130_fd_sc_hd__or2_1
XFILLER_47_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3985_ _5104_/Q _3983_/X _3980_/X _4833_/C vssd1 vssd1 vccd1 vccd1 _5104_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2936_ _2948_/A _2948_/B _2948_/C vssd1 vssd1 vccd1 vccd1 _2938_/A sky130_fd_sc_hd__nand3_1
X_2867_ _2863_/X _2864_/X _2865_/X _2866_/X vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__a22o_1
XFILLER_136_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4606_ _4606_/A vssd1 vssd1 vccd1 vccd1 _5304_/D sky130_fd_sc_hd__clkbuf_1
X_2798_ _5129_/Q vssd1 vssd1 vccd1 vccd1 _2870_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5586_ _5586_/A _2615_/Y vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__ebufn_8
X_4537_ _5282_/Q _5429_/Q _4541_/S vssd1 vssd1 vccd1 vccd1 _4538_/A sky130_fd_sc_hd__mux2_1
X_4468_ _4468_/A vssd1 vssd1 vccd1 vccd1 _5255_/D sky130_fd_sc_hd__clkbuf_1
X_3419_ _4073_/D _3419_/B vssd1 vssd1 vccd1 vccd1 _3420_/S sky130_fd_sc_hd__nand2_4
X_4399_ _5200_/Q _5170_/Q _4399_/S vssd1 vssd1 vccd1 vccd1 _4400_/B sky130_fd_sc_hd__mux2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3770_ _3741_/X _3768_/Y _3769_/X _3606_/A vssd1 vssd1 vccd1 vccd1 _3770_/X sky130_fd_sc_hd__a22o_1
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2721_ _2782_/A _2780_/A _2721_/C vssd1 vssd1 vccd1 vccd1 _2727_/A sky130_fd_sc_hd__and3_4
XFILLER_13_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5440_ _5443_/CLK _5440_/D vssd1 vssd1 vccd1 vccd1 _5440_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_9_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2652_ _2653_/A vssd1 vssd1 vccd1 vccd1 _2652_/Y sky130_fd_sc_hd__inv_2
X_2583_ _2585_/A vssd1 vssd1 vccd1 vccd1 _2583_/Y sky130_fd_sc_hd__inv_2
X_5371_ _5371_/CLK _5371_/D vssd1 vssd1 vccd1 vccd1 _5561_/A sky130_fd_sc_hd__dfxtp_1
X_4322_ _4322_/A vssd1 vssd1 vccd1 vccd1 _5221_/D sky130_fd_sc_hd__clkbuf_1
X_4253_ _4253_/A vssd1 vssd1 vccd1 vccd1 _5204_/D sky130_fd_sc_hd__clkbuf_1
X_5498__88 vssd1 vssd1 vccd1 vccd1 _5498__88/HI _5597_/A sky130_fd_sc_hd__conb_1
X_3204_ _5058_/Q vssd1 vssd1 vccd1 vccd1 _3424_/A sky130_fd_sc_hd__clkbuf_1
X_4184_ _4182_/X _5184_/Q _4197_/S vssd1 vssd1 vccd1 vccd1 _4185_/A sky130_fd_sc_hd__mux2_1
X_3135_ _3135_/A _3135_/B vssd1 vssd1 vccd1 vccd1 _4833_/C sky130_fd_sc_hd__xnor2_4
X_3066_ _3056_/X _3066_/B _3066_/C vssd1 vssd1 vccd1 vccd1 _3067_/C sky130_fd_sc_hd__nand3b_1
XFILLER_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3968_ _4906_/A vssd1 vssd1 vccd1 vccd1 _5437_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2919_ _2977_/A _2918_/X _5233_/Q vssd1 vssd1 vccd1 vccd1 _2919_/X sky130_fd_sc_hd__mux2_1
X_3899_ _4827_/A _3899_/B vssd1 vssd1 vccd1 vccd1 _3959_/S sky130_fd_sc_hd__and2_2
XFILLER_136_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5638_ _5638_/A _2677_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[34] sky130_fd_sc_hd__ebufn_8
X_5569_ _5569_/A _2594_/Y vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__ebufn_8
Xhold140 _5177_/Q vssd1 vssd1 vccd1 vccd1 _4161_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_46_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4940_ _5435_/Q _2889_/A _4940_/S vssd1 vssd1 vccd1 vccd1 _4941_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4871_ _5378_/D _4863_/X _4870_/Y _4861_/X vssd1 vssd1 vccd1 vccd1 _5410_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1_0__1652_ clkbuf_0__1652_/X vssd1 vssd1 vccd1 vccd1 _3996__4/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3822_ _3829_/B _3829_/C vssd1 vssd1 vccd1 vccd1 _3828_/A sky130_fd_sc_hd__and2_1
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3753_ _3753_/A0 _3753_/A1 _3773_/S vssd1 vssd1 vccd1 vccd1 _3753_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3684_ _5008_/Q _4266_/S _3682_/X hold134/X vssd1 vssd1 vccd1 vccd1 _5008_/D sky130_fd_sc_hd__a22o_1
X_2704_ _5046_/Q _5045_/Q _5048_/Q _5047_/Q vssd1 vssd1 vccd1 vccd1 _2705_/D sky130_fd_sc_hd__or4_1
X_2635_ _2635_/A vssd1 vssd1 vccd1 vccd1 _2640_/A sky130_fd_sc_hd__clkbuf_4
X_5423_ _5430_/CLK _5423_/D vssd1 vssd1 vccd1 vccd1 _5423_/Q sky130_fd_sc_hd__dfxtp_1
X_5354_ _5446_/CLK _5354_/D vssd1 vssd1 vccd1 vccd1 _5354_/Q sky130_fd_sc_hd__dfxtp_1
X_2566_ _2690_/A vssd1 vssd1 vccd1 vccd1 _2698_/A sky130_fd_sc_hd__buf_6
X_4305_ _4304_/X _5217_/Q _4309_/S vssd1 vssd1 vccd1 vccd1 _4306_/A sky130_fd_sc_hd__mux2_1
X_5285_ _5435_/CLK _5285_/D vssd1 vssd1 vccd1 vccd1 _5285_/Q sky130_fd_sc_hd__dfxtp_1
X_4236_ _4236_/A vssd1 vssd1 vccd1 vccd1 _5199_/D sky130_fd_sc_hd__clkbuf_1
X_4167_ _5179_/Q _4164_/A _4165_/Y vssd1 vssd1 vccd1 vccd1 _4167_/Y sky130_fd_sc_hd__o21bai_1
X_3118_ _3146_/A _3117_/Y _3118_/S vssd1 vssd1 vccd1 vccd1 _3119_/B sky130_fd_sc_hd__mux2_2
XFILLER_28_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4098_ hold88/A _4101_/C vssd1 vssd1 vccd1 vccd1 _4100_/A sky130_fd_sc_hd__and2_1
XFILLER_28_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3049_ _3108_/A _3051_/A _5394_/Q vssd1 vssd1 vccd1 vccd1 _3057_/A sky130_fd_sc_hd__and3_1
XFILLER_24_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5070_ _5077_/CLK _5070_/D vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
X_5468__58 vssd1 vssd1 vccd1 vccd1 _5468__58/HI _5545_/A sky130_fd_sc_hd__conb_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4021_ _4827_/A _5120_/Q vssd1 vssd1 vccd1 vccd1 _4022_/B sky130_fd_sc_hd__and2_1
XFILLER_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4923_ _5427_/Q _5378_/Q _4927_/S vssd1 vssd1 vccd1 vccd1 _4924_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4854_ _5407_/Q _4855_/B vssd1 vssd1 vccd1 vccd1 _4864_/C sky130_fd_sc_hd__and2_1
X_4785_ _4785_/A _4785_/B vssd1 vssd1 vccd1 vccd1 _5368_/D sky130_fd_sc_hd__nor2_1
X_3805_ _3810_/C _3805_/B _3805_/C vssd1 vssd1 vccd1 vccd1 _3806_/A sky130_fd_sc_hd__and3b_1
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3736_ _3736_/A vssd1 vssd1 vccd1 vccd1 _3736_/Y sky130_fd_sc_hd__inv_2
X_3667_ _3667_/A _3667_/B vssd1 vssd1 vccd1 vccd1 _4276_/A sky130_fd_sc_hd__nor2_2
X_5406_ _5403_/Q _5406_/D vssd1 vssd1 vccd1 vccd1 _5406_/Q sky130_fd_sc_hd__dfxtp_1
X_2618_ _2622_/A vssd1 vssd1 vccd1 vccd1 _2618_/Y sky130_fd_sc_hd__inv_2
X_3598_ _3705_/A _3705_/B _3705_/C _3705_/D vssd1 vssd1 vccd1 vccd1 _3750_/B sky130_fd_sc_hd__or4_2
X_2549_ _2549_/A vssd1 vssd1 vccd1 vccd1 _5116_/D sky130_fd_sc_hd__clkbuf_1
X_5337_ _5446_/CLK _5337_/D vssd1 vssd1 vccd1 vccd1 _5337_/Q sky130_fd_sc_hd__dfxtp_1
X_5268_ _5322_/CLK _5268_/D vssd1 vssd1 vccd1 vccd1 _5268_/Q sky130_fd_sc_hd__dfxtp_1
X_4219_ _4611_/A vssd1 vssd1 vccd1 vccd1 _4235_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5199_ _5369_/CLK _5199_/D vssd1 vssd1 vccd1 vccd1 _5199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5482__72 vssd1 vssd1 vccd1 vccd1 _5482__72/HI _5559_/A sky130_fd_sc_hd__conb_1
XFILLER_51_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4570_ _5295_/Q _4577_/B vssd1 vssd1 vccd1 vccd1 _4570_/X sky130_fd_sc_hd__or2_1
XFILLER_7_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3521_ _4434_/A _3511_/Y _4220_/C _3658_/A vssd1 vssd1 vccd1 vccd1 _3524_/A sky130_fd_sc_hd__a211oi_1
X_3452_ _3476_/A _2874_/X _2875_/X _3476_/B vssd1 vssd1 vccd1 vccd1 _3452_/X sky130_fd_sc_hd__a22o_1
X_3383_ _3350_/S _3267_/A _3357_/X _3268_/A vssd1 vssd1 vccd1 vccd1 _3383_/X sky130_fd_sc_hd__o211a_1
X_5122_ _5439_/CLK _5122_/D vssd1 vssd1 vccd1 vccd1 _5586_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_57_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5053_ _5064_/CLK _5053_/D vssd1 vssd1 vccd1 vccd1 _5053_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _4906_/A _5436_/D vssd1 vssd1 vccd1 vccd1 _4940_/S sky130_fd_sc_hd__or2_2
XFILLER_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4837_ _5230_/Q _4837_/B vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__and2b_1
X_4768_ _5363_/Q _4771_/C vssd1 vssd1 vccd1 vccd1 _4774_/C sky130_fd_sc_hd__and2_1
X_4699_ _4589_/Y _4698_/X _4588_/X vssd1 vssd1 vccd1 vccd1 _4700_/C sky130_fd_sc_hd__o21ai_1
X_3719_ _4022_/A vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__clkbuf_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__clkbuf_2
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_8 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2952_ _2953_/B _2977_/C vssd1 vssd1 vccd1 vccd1 _2952_/Y sky130_fd_sc_hd__nor2_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2883_ _5239_/Q vssd1 vssd1 vccd1 vccd1 _2950_/A sky130_fd_sc_hd__inv_2
X_4622_ _4666_/S vssd1 vssd1 vccd1 vccd1 _4640_/S sky130_fd_sc_hd__buf_2
X_4553_ _4553_/A _4587_/C _4594_/B vssd1 vssd1 vccd1 vccd1 _4581_/B sky130_fd_sc_hd__and3_1
X_4484_ _5262_/Q _5100_/Q _4492_/S vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__mux2_1
X_3504_ _4112_/A _3673_/B vssd1 vssd1 vccd1 vccd1 _3528_/A sky130_fd_sc_hd__nor2_1
X_3435_ _5134_/Q vssd1 vssd1 vccd1 vccd1 _5629_/A sky130_fd_sc_hd__clkinv_2
X_3366_ _3361_/X _3363_/X _3373_/B vssd1 vssd1 vccd1 vccd1 _3366_/Y sky130_fd_sc_hd__a21oi_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3297_ _4995_/Q _3295_/B _4996_/Q vssd1 vssd1 vccd1 vccd1 _3553_/A sky130_fd_sc_hd__o21ai_2
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5437_/CLK _5105_/D vssd1 vssd1 vccd1 vccd1 _5105_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5439_/CLK _5036_/D vssd1 vssd1 vccd1 vccd1 _5036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3220_ _3445_/C _3191_/A _5440_/Q vssd1 vssd1 vccd1 vccd1 _3221_/C sky130_fd_sc_hd__a21o_1
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3151_ _3150_/A _3150_/B _3150_/C vssd1 vssd1 vccd1 vccd1 _3166_/B sky130_fd_sc_hd__a21o_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3082_ _3081_/A _3081_/B _3081_/C vssd1 vssd1 vccd1 vccd1 _3102_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3984_ _5103_/Q _3983_/X _3980_/X _4834_/B vssd1 vssd1 vccd1 vccd1 _5103_/D sky130_fd_sc_hd__a22o_1
X_2935_ _2934_/B _2934_/C _5236_/Q vssd1 vssd1 vccd1 vccd1 _2948_/C sky130_fd_sc_hd__a21o_1
X_2866_ _2870_/B _2870_/A vssd1 vssd1 vccd1 vccd1 _2866_/X sky130_fd_sc_hd__and2b_1
XFILLER_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4605_ _4609_/A _4605_/B vssd1 vssd1 vccd1 vccd1 _4606_/A sky130_fd_sc_hd__and2_1
X_2797_ _2840_/A vssd1 vssd1 vccd1 vccd1 _2870_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5585_ _5585_/A _2614_/Y vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__ebufn_8
X_4536_ _4536_/A vssd1 vssd1 vccd1 vccd1 _5281_/D sky130_fd_sc_hd__clkbuf_1
X_4467_ _5255_/Q _5093_/Q _4583_/B vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__mux2_1
X_3418_ _5126_/Q _5125_/Q _3418_/S vssd1 vssd1 vccd1 vccd1 _3418_/X sky130_fd_sc_hd__mux2_1
X_4398_ _3652_/A _4383_/X _4396_/X _4397_/X vssd1 vssd1 vccd1 vccd1 _5236_/D sky130_fd_sc_hd__o211a_1
X_3349_ _3349_/A _3349_/B vssd1 vssd1 vccd1 vccd1 _3350_/S sky130_fd_sc_hd__nand2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5518__108 vssd1 vssd1 vccd1 vccd1 _5518__108/HI _5634_/A sky130_fd_sc_hd__conb_1
X_5019_ _5058_/CLK _5019_/D vssd1 vssd1 vccd1 vccd1 _5019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2720_ _2717_/X _2778_/A _2720_/C vssd1 vssd1 vccd1 vccd1 _2721_/C sky130_fd_sc_hd__and3b_1
XFILLER_13_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2651_ _2653_/A vssd1 vssd1 vccd1 vccd1 _2651_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2582_ _2585_/A vssd1 vssd1 vccd1 vccd1 _2582_/Y sky130_fd_sc_hd__inv_2
X_5370_ _5446_/CLK _5370_/D vssd1 vssd1 vccd1 vccd1 _5370_/Q sky130_fd_sc_hd__dfxtp_1
X_4321_ _4320_/X _5221_/Q _4324_/S vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__mux2_1
XFILLER_4_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4252_ _4252_/A _4252_/B vssd1 vssd1 vccd1 vccd1 _4253_/A sky130_fd_sc_hd__and2_1
X_3203_ _5052_/Q vssd1 vssd1 vccd1 vccd1 _3823_/D sky130_fd_sc_hd__inv_2
X_4183_ _4200_/A vssd1 vssd1 vccd1 vccd1 _4197_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3134_ _3134_/A _3134_/B vssd1 vssd1 vccd1 vccd1 _3135_/B sky130_fd_sc_hd__xnor2_2
X_3065_ _3065_/A vssd1 vssd1 vccd1 vccd1 _3067_/A sky130_fd_sc_hd__clkinv_2
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3967_ _3967_/A _4904_/C vssd1 vssd1 vccd1 vccd1 _4906_/A sky130_fd_sc_hd__nor2_1
X_2918_ _4831_/A vssd1 vssd1 vccd1 vccd1 _2918_/X sky130_fd_sc_hd__clkbuf_4
X_3898_ _5278_/Q _3910_/A _3897_/X _5014_/Q vssd1 vssd1 vccd1 vccd1 _3898_/X sky130_fd_sc_hd__a22o_1
X_5637_ _5637_/A _2676_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[33] sky130_fd_sc_hd__ebufn_8
X_2849_ _2825_/Y _2837_/X _2848_/X _2817_/S vssd1 vssd1 vccd1 vccd1 _2849_/X sky130_fd_sc_hd__a22o_1
X_5568_ _5568_/A _2593_/Y vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__ebufn_8
Xhold130 _5062_/Q vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold141 _5274_/Q vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_4519_ _5274_/Q _5421_/Q _4519_/S vssd1 vssd1 vccd1 vccd1 _4520_/A sky130_fd_sc_hd__mux2_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4870_ _4875_/C _4869_/Y _4851_/X vssd1 vssd1 vccd1 vccd1 _4870_/Y sky130_fd_sc_hd__o21ai_1
X_3821_ _3821_/A vssd1 vssd1 vccd1 vccd1 _5051_/D sky130_fd_sc_hd__clkbuf_1
X_3752_ _3752_/A vssd1 vssd1 vccd1 vccd1 _3773_/S sky130_fd_sc_hd__buf_2
X_3683_ _5007_/Q _4266_/S _3682_/X hold142/X vssd1 vssd1 vccd1 vccd1 _5007_/D sky130_fd_sc_hd__a22o_1
X_2703_ _5042_/Q _5041_/Q _5044_/Q _5043_/Q vssd1 vssd1 vccd1 vccd1 _2706_/A sky130_fd_sc_hd__or4_1
X_2634_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2634_/Y sky130_fd_sc_hd__inv_2
X_5422_ _5430_/CLK _5422_/D vssd1 vssd1 vccd1 vccd1 _5422_/Q sky130_fd_sc_hd__dfxtp_1
X_2565_ input1/X vssd1 vssd1 vccd1 vccd1 _2690_/A sky130_fd_sc_hd__buf_6
X_5353_ _5353_/CLK _5353_/D vssd1 vssd1 vccd1 vccd1 _5353_/Q sky130_fd_sc_hd__dfxtp_1
X_4304_ _5213_/Q _4264_/X _4303_/X vssd1 vssd1 vccd1 vccd1 _4304_/X sky130_fd_sc_hd__a21o_1
X_5284_ _5431_/CLK _5284_/D vssd1 vssd1 vccd1 vccd1 _5284_/Q sky130_fd_sc_hd__dfxtp_1
X_4235_ _4235_/A _4235_/B vssd1 vssd1 vccd1 vccd1 _4236_/A sky130_fd_sc_hd__and2_1
X_4166_ _5178_/Q _4163_/B _4164_/Y _4165_/Y vssd1 vssd1 vccd1 vccd1 _5178_/D sky130_fd_sc_hd__a211o_1
X_3117_ _3144_/B _3117_/B vssd1 vssd1 vccd1 vccd1 _3117_/Y sky130_fd_sc_hd__xnor2_1
X_4097_ _2727_/A _5148_/Q vssd1 vssd1 vccd1 vccd1 _4101_/C sky130_fd_sc_hd__and2b_1
X_3048_ _3040_/A _3040_/B _3041_/A _3036_/A vssd1 vssd1 vccd1 vccd1 _3060_/A sky130_fd_sc_hd__o211ai_4
XFILLER_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4999_ _5058_/CLK _4999_/D vssd1 vssd1 vccd1 vccd1 _4999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_17_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5323_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4020_ _4020_/A vssd1 vssd1 vccd1 vccd1 _5126_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4922_ _4922_/A vssd1 vssd1 vccd1 vccd1 _5426_/D sky130_fd_sc_hd__clkbuf_1
X_4853_ _5374_/D _4840_/X _4852_/Y _4842_/X vssd1 vssd1 vccd1 vccd1 _5406_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4784_ _5368_/Q _4782_/A _4742_/X vssd1 vssd1 vccd1 vccd1 _4785_/B sky130_fd_sc_hd__o21ai_1
X_3804_ _5044_/Q _5045_/Q _3797_/B _5046_/Q vssd1 vssd1 vccd1 vccd1 _3805_/B sky130_fd_sc_hd__a31o_1
X_3735_ _5022_/Q _3767_/A _3731_/Y _3734_/X vssd1 vssd1 vccd1 vccd1 _5022_/D sky130_fd_sc_hd__a211o_1
X_5405_ _5403_/Q _5405_/D vssd1 vssd1 vccd1 vccd1 _5405_/Q sky130_fd_sc_hd__dfxtp_1
X_3666_ _4112_/A _4434_/C vssd1 vssd1 vccd1 vccd1 _3667_/B sky130_fd_sc_hd__nand2_1
X_2617_ _2635_/A vssd1 vssd1 vccd1 vccd1 _2622_/A sky130_fd_sc_hd__clkbuf_2
X_3597_ _5040_/Q _2753_/B _3715_/A vssd1 vssd1 vccd1 vccd1 _3597_/X sky130_fd_sc_hd__o21a_1
X_2548_ _2541_/B _2548_/B _2548_/C vssd1 vssd1 vccd1 vccd1 _2549_/A sky130_fd_sc_hd__and3b_1
X_5336_ _5446_/CLK _5336_/D vssd1 vssd1 vccd1 vccd1 _5336_/Q sky130_fd_sc_hd__dfxtp_1
X_5267_ _5328_/CLK _5267_/D vssd1 vssd1 vccd1 vccd1 _5267_/Q sky130_fd_sc_hd__dfxtp_1
X_4218_ _4218_/A vssd1 vssd1 vccd1 vccd1 _5194_/D sky130_fd_sc_hd__clkbuf_1
X_5198_ _5369_/CLK _5198_/D vssd1 vssd1 vccd1 vccd1 _5198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4149_ _4149_/A vssd1 vssd1 vccd1 vccd1 _5175_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3520_ _3531_/A _3519_/X _4355_/C vssd1 vssd1 vccd1 vccd1 _3658_/A sky130_fd_sc_hd__o21ai_1
XFILLER_7_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3451_ _2864_/X _2865_/X _3450_/X vssd1 vssd1 vccd1 vccd1 _3451_/Y sky130_fd_sc_hd__a21oi_1
X_3382_ _3352_/S _3267_/X _3378_/Y _3381_/X vssd1 vssd1 vccd1 vccd1 _3382_/X sky130_fd_sc_hd__a31o_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5121_ _5121_/CLK _5121_/D vssd1 vssd1 vccd1 vccd1 _5121_/Q sky130_fd_sc_hd__dfxtp_1
X_5052_ _5439_/CLK _5052_/D vssd1 vssd1 vccd1 vccd1 _5052_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4905_ _4905_/A vssd1 vssd1 vccd1 vccd1 _5436_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4836_ _3170_/X _3186_/X _4835_/C _5228_/Q vssd1 vssd1 vccd1 vccd1 _4836_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4767_ _4771_/C _4767_/B vssd1 vssd1 vccd1 vccd1 _5362_/D sky130_fd_sc_hd__nor2_1
X_3718_ _3718_/A _3724_/B vssd1 vssd1 vccd1 vccd1 _3718_/Y sky130_fd_sc_hd__nand2_1
X_4698_ _5327_/Q _4698_/B vssd1 vssd1 vccd1 vccd1 _4698_/X sky130_fd_sc_hd__and2_1
X_3649_ _3649_/A _3649_/B vssd1 vssd1 vccd1 vccd1 _3649_/Y sky130_fd_sc_hd__nand2_1
X_5319_ _5322_/CLK _5319_/D vssd1 vssd1 vccd1 vccd1 _5574_/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_9 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2951_ _5238_/Q _2951_/B vssd1 vssd1 vccd1 vccd1 _2962_/A sky130_fd_sc_hd__xnor2_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2882_ _2953_/B vssd1 vssd1 vccd1 vccd1 _2977_/A sky130_fd_sc_hd__clkbuf_4
X_4621_ _5290_/Q _5260_/Q _4639_/S vssd1 vssd1 vccd1 vccd1 _4621_/X sky130_fd_sc_hd__mux2_1
X_4552_ _4566_/A vssd1 vssd1 vccd1 vccd1 _4552_/X sky130_fd_sc_hd__clkbuf_2
X_4483_ _4532_/A vssd1 vssd1 vccd1 vccd1 _4492_/S sky130_fd_sc_hd__clkbuf_2
X_3503_ _5247_/Q vssd1 vssd1 vccd1 vccd1 _3673_/B sky130_fd_sc_hd__inv_2
X_3434_ _5245_/Q vssd1 vssd1 vccd1 vccd1 _5623_/A sky130_fd_sc_hd__clkinv_4
X_3365_ _3344_/A _3364_/Y _3338_/A vssd1 vssd1 vccd1 vccd1 _3373_/B sky130_fd_sc_hd__o21a_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3296_ _3396_/A _3305_/B _3302_/A vssd1 vssd1 vccd1 vccd1 _3298_/A sky130_fd_sc_hd__o21a_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _5436_/CLK _5104_/D vssd1 vssd1 vccd1 vccd1 _5104_/Q sky130_fd_sc_hd__dfxtp_1
X_5035_ _5058_/CLK _5035_/D vssd1 vssd1 vccd1 vccd1 _5035_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3995__3 _3996__4/A vssd1 vssd1 vccd1 vccd1 _5110_/CLK sky130_fd_sc_hd__inv_2
XFILLER_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4819_ _4834_/C _5399_/Q _4823_/S vssd1 vssd1 vccd1 vccd1 _4820_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3150_ _3150_/A _3150_/B _3150_/C vssd1 vssd1 vccd1 vccd1 _3152_/A sky130_fd_sc_hd__and3_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3081_ _3081_/A _3081_/B _3081_/C vssd1 vssd1 vccd1 vccd1 _3081_/Y sky130_fd_sc_hd__nand3_1
XFILLER_35_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3983_ _3983_/A vssd1 vssd1 vccd1 vccd1 _3983_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2934_ _5236_/Q _2934_/B _2934_/C vssd1 vssd1 vccd1 vccd1 _2948_/B sky130_fd_sc_hd__nand3_1
X_2865_ _4998_/Q _5035_/Q _2869_/A vssd1 vssd1 vccd1 vccd1 _2865_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4604_ _5304_/Q _4603_/X _4617_/S vssd1 vssd1 vccd1 vccd1 _4605_/B sky130_fd_sc_hd__mux2_1
X_5584_ _5584_/A _2613_/Y vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__ebufn_8
X_2796_ _5128_/Q vssd1 vssd1 vccd1 vccd1 _2840_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4535_ _5281_/Q _5428_/Q _4541_/S vssd1 vssd1 vccd1 vccd1 _4536_/A sky130_fd_sc_hd__mux2_1
X_4466_ _4532_/A vssd1 vssd1 vccd1 vccd1 _4583_/B sky130_fd_sc_hd__clkbuf_2
X_3417_ _5124_/Q _5123_/Q _3418_/S vssd1 vssd1 vccd1 vccd1 _3417_/X sky130_fd_sc_hd__mux2_1
X_4397_ _4667_/A vssd1 vssd1 vccd1 vccd1 _4397_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3348_ _3563_/A _3419_/B vssd1 vssd1 vccd1 vccd1 _3348_/X sky130_fd_sc_hd__and2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3279_ _5443_/Q _3279_/B vssd1 vssd1 vccd1 vccd1 _3279_/Y sky130_fd_sc_hd__xnor2_1
X_5018_ _5058_/CLK _5018_/D vssd1 vssd1 vccd1 vccd1 _5018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2650_ _2653_/A vssd1 vssd1 vccd1 vccd1 _2650_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2581_ _2585_/A vssd1 vssd1 vccd1 vccd1 _2581_/Y sky130_fd_sc_hd__inv_2
X_4320_ _5217_/Q _3535_/X _3537_/X _5171_/Q _3543_/B vssd1 vssd1 vccd1 vccd1 _4320_/X
+ sky130_fd_sc_hd__a221o_1
X_4251_ _5204_/Q _5200_/Q _4251_/S vssd1 vssd1 vccd1 vccd1 _4252_/B sky130_fd_sc_hd__mux2_1
X_3202_ _3216_/A vssd1 vssd1 vccd1 vccd1 _3829_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4182_ _5408_/Q _5359_/Q _4182_/S vssd1 vssd1 vccd1 vccd1 _4182_/X sky130_fd_sc_hd__mux2_1
X_3133_ _3084_/A _3146_/B _3132_/X vssd1 vssd1 vccd1 vccd1 _3134_/B sky130_fd_sc_hd__a21bo_1
X_3064_ _5379_/Q _3028_/X _4832_/C _3009_/X _3063_/X vssd1 vssd1 vccd1 vccd1 _5379_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3966_ _3983_/A vssd1 vssd1 vccd1 vccd1 _3966_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2917_ _2939_/A _2917_/B vssd1 vssd1 vccd1 vccd1 _4831_/A sky130_fd_sc_hd__xnor2_1
X_5636_ _5636_/A _2675_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[32] sky130_fd_sc_hd__ebufn_8
X_3897_ _3903_/A vssd1 vssd1 vccd1 vccd1 _3897_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2848_ _2838_/X _2843_/X _2847_/X _2825_/Y vssd1 vssd1 vccd1 vccd1 _2848_/X sky130_fd_sc_hd__a22o_1
X_5567_ _5567_/A _2591_/Y vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__ebufn_8
X_2779_ _5153_/Q _5152_/Q _5151_/Q vssd1 vssd1 vccd1 vccd1 _2781_/B sky130_fd_sc_hd__and3_1
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__clkbuf_1
Xhold142 _5183_/Q vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_4518_ _5273_/Q _4512_/A _4517_/Y vssd1 vssd1 vccd1 vccd1 _5273_/D sky130_fd_sc_hd__a21o_1
X_4449_ _5251_/Q _4449_/B _4449_/C vssd1 vssd1 vccd1 vccd1 _4455_/B sky130_fd_sc_hd__and3_1
X_5489__79 vssd1 vssd1 vccd1 vccd1 _5489__79/HI _5567_/A sky130_fd_sc_hd__conb_1
XFILLER_58_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _3820_/A _3820_/B _3820_/C vssd1 vssd1 vccd1 vccd1 _3821_/A sky130_fd_sc_hd__and3_1
X_3751_ _3751_/A _3751_/B vssd1 vssd1 vccd1 vccd1 _3751_/Y sky130_fd_sc_hd__nand2_1
X_2702_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4348_/A sky130_fd_sc_hd__clkbuf_4
X_3682_ _4350_/A _3682_/B _3682_/C _3682_/D vssd1 vssd1 vccd1 vccd1 _3682_/X sky130_fd_sc_hd__and4_2
X_2633_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2633_/Y sky130_fd_sc_hd__inv_2
X_5421_ _5430_/CLK _5421_/D vssd1 vssd1 vccd1 vccd1 _5421_/Q sky130_fd_sc_hd__dfxtp_1
X_5352_ _5353_/CLK _5352_/D vssd1 vssd1 vccd1 vccd1 _5352_/Q sky130_fd_sc_hd__dfxtp_1
X_2564_ _2564_/A _2564_/B vssd1 vssd1 vccd1 vccd1 _5110_/D sky130_fd_sc_hd__nor2_1
X_4303_ _5167_/Q _4285_/X _4276_/A _5193_/Q vssd1 vssd1 vccd1 vccd1 _4303_/X sky130_fd_sc_hd__a22o_1
X_5283_ _5431_/CLK _5283_/D vssd1 vssd1 vccd1 vccd1 _5283_/Q sky130_fd_sc_hd__dfxtp_1
X_4234_ _5199_/Q _5195_/Q _4234_/S vssd1 vssd1 vccd1 vccd1 _4235_/B sky130_fd_sc_hd__mux2_1
X_4165_ _4165_/A _4165_/B vssd1 vssd1 vccd1 vccd1 _4165_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3116_ _3102_/B _3115_/X _3099_/A vssd1 vssd1 vccd1 vccd1 _3117_/B sky130_fd_sc_hd__a21o_1
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4096_ _5155_/Q _4093_/C _4095_/Y vssd1 vssd1 vccd1 vccd1 _5155_/D sky130_fd_sc_hd__o21a_1
X_3047_ _5378_/Q _3028_/X _4833_/A _3009_/X _3046_/X vssd1 vssd1 vccd1 vccd1 _5378_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_36_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4998_ _5058_/CLK _4998_/D vssd1 vssd1 vccd1 vccd1 _4998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3949_ _5085_/Q _3943_/X _3948_/X _3911_/X vssd1 vssd1 vccd1 vccd1 _3949_/X sky130_fd_sc_hd__a211o_1
XFILLER_137_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5619_ _5619_/A _2655_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[15] sky130_fd_sc_hd__ebufn_8
XFILLER_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4921_ _5426_/Q _5377_/Q _4927_/S vssd1 vssd1 vccd1 vccd1 _4922_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4852_ _4849_/Y _4855_/B _4851_/X vssd1 vssd1 vccd1 vccd1 _4852_/Y sky130_fd_sc_hd__o21ai_1
X_3803_ _5046_/Q _5045_/Q _3803_/C vssd1 vssd1 vccd1 vccd1 _3810_/C sky130_fd_sc_hd__and3_1
XFILLER_21_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4783_ _5368_/Q _5367_/Q _4783_/C vssd1 vssd1 vccd1 vccd1 _4785_/A sky130_fd_sc_hd__and3_1
X_3734_ _3734_/A _3734_/B _3740_/A vssd1 vssd1 vccd1 vccd1 _3734_/X sky130_fd_sc_hd__and3_1
X_3665_ _3665_/A vssd1 vssd1 vccd1 vccd1 _4165_/A sky130_fd_sc_hd__clkbuf_2
X_5404_ _5403_/Q _5404_/D vssd1 vssd1 vccd1 vccd1 _5404_/Q sky130_fd_sc_hd__dfxtp_1
X_2616_ _2616_/A vssd1 vssd1 vccd1 vccd1 _2616_/Y sky130_fd_sc_hd__inv_2
X_3596_ _3596_/A _3720_/B vssd1 vssd1 vccd1 vccd1 _3604_/B sky130_fd_sc_hd__nor2_1
X_5335_ _5335_/CLK _5335_/D vssd1 vssd1 vccd1 vccd1 _5335_/Q sky130_fd_sc_hd__dfxtp_1
X_2547_ _2734_/A _2554_/A _5116_/Q vssd1 vssd1 vccd1 vccd1 _2548_/B sky130_fd_sc_hd__a21o_1
X_5459__49 vssd1 vssd1 vccd1 vccd1 _5459__49/HI _5536_/A sky130_fd_sc_hd__conb_1
X_5266_ _5322_/CLK _5266_/D vssd1 vssd1 vccd1 vccd1 _5266_/Q sky130_fd_sc_hd__dfxtp_1
X_4217_ _4216_/X _5194_/Q _4261_/S vssd1 vssd1 vccd1 vccd1 _4218_/A sky130_fd_sc_hd__mux2_1
X_5197_ _5445_/CLK _5197_/D vssd1 vssd1 vccd1 vccd1 _5197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4148_ _5352_/Q _5175_/Q _4148_/S vssd1 vssd1 vccd1 vccd1 _4149_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4079_ _4084_/B _4080_/A vssd1 vssd1 vccd1 vccd1 _4083_/A sky130_fd_sc_hd__and2_1
XFILLER_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5473__63 vssd1 vssd1 vccd1 vccd1 _5473__63/HI _5550_/A sky130_fd_sc_hd__conb_1
XFILLER_61_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3450_ _3476_/A _2863_/X _2868_/X _3476_/B vssd1 vssd1 vccd1 vccd1 _3450_/X sky130_fd_sc_hd__a22o_1
X_3381_ _3378_/B _3380_/B _3380_/Y _3357_/X vssd1 vssd1 vccd1 vccd1 _3381_/X sky130_fd_sc_hd__o22a_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5120_ _5120_/CLK _5120_/D vssd1 vssd1 vccd1 vccd1 _5120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5051_ _5051_/CLK _5051_/D vssd1 vssd1 vccd1 vccd1 _5051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4904_ _4829_/S _5419_/Q _4904_/C vssd1 vssd1 vccd1 vccd1 _4905_/A sky130_fd_sc_hd__and3b_1
XFILLER_21_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4835_ _4835_/A _4835_/B _4835_/C _5229_/Q vssd1 vssd1 vccd1 vccd1 _4835_/X sky130_fd_sc_hd__or4b_1
X_4766_ _5362_/Q _4764_/A _4762_/X vssd1 vssd1 vccd1 vccd1 _4767_/B sky130_fd_sc_hd__o21ai_1
X_3717_ _3729_/A _3734_/B _3754_/B vssd1 vssd1 vccd1 vccd1 _3724_/B sky130_fd_sc_hd__and3_1
X_4697_ _4587_/C _4693_/B _4698_/B _5327_/Q vssd1 vssd1 vccd1 vccd1 _4700_/B sky130_fd_sc_hd__a31o_1
XFILLER_136_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3648_ _3648_/A _3648_/B vssd1 vssd1 vccd1 vccd1 _3649_/B sky130_fd_sc_hd__xnor2_1
X_3579_ _4073_/C _3577_/A _3569_/X vssd1 vssd1 vccd1 vccd1 _3580_/B sky130_fd_sc_hd__o21ai_1
X_5318_ _5437_/CLK _5318_/D vssd1 vssd1 vccd1 vccd1 _5318_/Q sky130_fd_sc_hd__dfxtp_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _5446_/CLK _5249_/D vssd1 vssd1 vccd1 vccd1 _5249_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_2_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5439_/CLK
+ sky130_fd_sc_hd__clkbuf_16
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2950_ _2950_/A _5389_/Q vssd1 vssd1 vccd1 vccd1 _2951_/B sky130_fd_sc_hd__and2_1
X_2881_ _5372_/Q vssd1 vssd1 vccd1 vccd1 _2953_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4665_/S vssd1 vssd1 vccd1 vccd1 _4639_/S sky130_fd_sc_hd__clkbuf_2
X_4551_ _4693_/A _4551_/B vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__nand2_2
XFILLER_7_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4482_ _4482_/A vssd1 vssd1 vccd1 vccd1 _5261_/D sky130_fd_sc_hd__clkbuf_1
X_3502_ _4730_/A vssd1 vssd1 vccd1 vccd1 _4112_/A sky130_fd_sc_hd__clkbuf_2
X_3433_ _5320_/Q vssd1 vssd1 vccd1 vccd1 _5617_/A sky130_fd_sc_hd__clkinv_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _3418_/S _3380_/A vssd1 vssd1 vccd1 vccd1 _3364_/Y sky130_fd_sc_hd__nor2_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5436_/CLK _5103_/D vssd1 vssd1 vccd1 vccd1 _5103_/Q sky130_fd_sc_hd__dfxtp_1
X_3295_ _4995_/Q _3295_/B vssd1 vssd1 vccd1 vccd1 _3302_/A sky130_fd_sc_hd__xnor2_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5058_/CLK _5034_/D vssd1 vssd1 vccd1 vccd1 _5034_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4818_ _4818_/A vssd1 vssd1 vccd1 vccd1 _5398_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4749_ _5357_/Q _4752_/C vssd1 vssd1 vccd1 vccd1 _4751_/A sky130_fd_sc_hd__and2_1
XFILLER_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3080_ _3083_/A _3083_/B vssd1 vssd1 vccd1 vccd1 _3081_/C sky130_fd_sc_hd__xnor2_1
XFILLER_47_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3982_ _5102_/Q _3976_/X _3980_/X _4834_/A vssd1 vssd1 vccd1 vccd1 _5102_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2933_ _5240_/Q _2902_/X _2910_/A vssd1 vssd1 vccd1 vccd1 _2934_/C sky130_fd_sc_hd__o21a_1
X_2864_ _2870_/A _2870_/B vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__and2b_1
X_2795_ _2833_/A vssd1 vssd1 vccd1 vccd1 _2795_/X sky130_fd_sc_hd__buf_2
X_4603_ input3/X _5256_/Q _4616_/S vssd1 vssd1 vccd1 vccd1 _4603_/X sky130_fd_sc_hd__mux2_1
X_5583_ _5583_/A _2612_/Y vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__ebufn_8
X_4534_ _4534_/A vssd1 vssd1 vccd1 vccd1 _5280_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4465_ _4471_/A vssd1 vssd1 vccd1 vccd1 _4532_/A sky130_fd_sc_hd__clkbuf_2
X_3416_ _3389_/Y _3395_/X _3414_/X _4902_/A vssd1 vssd1 vccd1 vccd1 _3416_/X sky130_fd_sc_hd__a31o_1
X_4396_ _4400_/A _4396_/B vssd1 vssd1 vccd1 vccd1 _4396_/X sky130_fd_sc_hd__or2_1
X_3347_ _4990_/Q vssd1 vssd1 vccd1 vccd1 _3563_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _5058_/CLK _5017_/D vssd1 vssd1 vccd1 vccd1 _5017_/Q sky130_fd_sc_hd__dfxtp_1
X_3278_ _3424_/C _3277_/Y _3285_/B vssd1 vssd1 vccd1 vccd1 _3279_/B sky130_fd_sc_hd__mux2_1
XFILLER_54_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2580_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2585_/A sky130_fd_sc_hd__buf_2
X_4250_ _4250_/A vssd1 vssd1 vccd1 vccd1 _5203_/D sky130_fd_sc_hd__clkbuf_1
X_3201_ _3285_/B _3229_/B vssd1 vssd1 vccd1 vccd1 _3275_/A sky130_fd_sc_hd__nand2_1
X_4181_ _4181_/A vssd1 vssd1 vccd1 vccd1 _5183_/D sky130_fd_sc_hd__clkbuf_1
X_3132_ _3132_/A _3132_/B _3132_/C vssd1 vssd1 vccd1 vccd1 _3132_/X sky130_fd_sc_hd__or3_1
XFILLER_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3063_ _3106_/A _3649_/A vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__or2_1
XFILLER_48_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3965_ _4829_/S _3961_/Y _4904_/C vssd1 vssd1 vccd1 vccd1 _3983_/A sky130_fd_sc_hd__o21a_2
XFILLER_50_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2916_ _5234_/Q _2916_/B vssd1 vssd1 vccd1 vccd1 _2917_/B sky130_fd_sc_hd__xnor2_1
X_3896_ _4692_/C _3946_/A _3945_/B _3942_/B vssd1 vssd1 vccd1 vccd1 _3903_/A sky130_fd_sc_hd__a31o_1
X_5635_ _5635_/A _2674_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__ebufn_8
X_2847_ _2844_/X _5032_/Q _5031_/Q _5034_/Q _2833_/X _2846_/X vssd1 vssd1 vccd1 vccd1
+ _2847_/X sky130_fd_sc_hd__mux4_1
XFILLER_12_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5566_ _5566_/A _2698_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__ebufn_8
X_2778_ _2778_/A _2778_/B vssd1 vssd1 vccd1 vccd1 _2785_/A sky130_fd_sc_hd__nor2_1
Xhold110 _5154_/Q vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold132 _5151_/Q vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold121 _5152_/Q vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_2_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold143 _5084_/Q vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_4517_ _5273_/Q _4512_/A _4515_/C vssd1 vssd1 vccd1 vccd1 _4517_/Y sky130_fd_sc_hd__o21bai_1
X_5524__114 vssd1 vssd1 vccd1 vccd1 _5524__114/HI _5640_/A sky130_fd_sc_hd__conb_1
X_4448_ _4445_/X _4446_/X _4447_/Y _4954_/A vssd1 vssd1 vccd1 vccd1 _5250_/D sky130_fd_sc_hd__a211oi_1
X_4379_ _5231_/Q _4362_/X _4376_/X _4378_/X vssd1 vssd1 vccd1 vccd1 _5231_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3750_ _3750_/A _3750_/B vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__and2_1
XFILLER_20_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2701_ _4708_/A vssd1 vssd1 vccd1 vccd1 _4094_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3681_ _3698_/A vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__buf_4
X_2632_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2632_/Y sky130_fd_sc_hd__inv_2
X_5420_ _5430_/CLK _5420_/D vssd1 vssd1 vccd1 vccd1 _5420_/Q sky130_fd_sc_hd__dfxtp_1
X_5351_ _5351_/CLK _5351_/D vssd1 vssd1 vccd1 vccd1 _5351_/Q sky130_fd_sc_hd__dfxtp_1
X_2563_ _3705_/C _2560_/B _2530_/B vssd1 vssd1 vccd1 vccd1 _2564_/B sky130_fd_sc_hd__o21ai_1
X_5282_ _5430_/CLK _5282_/D vssd1 vssd1 vccd1 vccd1 _5282_/Q sky130_fd_sc_hd__dfxtp_1
X_4302_ _4302_/A vssd1 vssd1 vccd1 vccd1 _5216_/D sky130_fd_sc_hd__clkbuf_1
X_4233_ _4233_/A vssd1 vssd1 vccd1 vccd1 _5198_/D sky130_fd_sc_hd__clkbuf_1
X_4164_ _4164_/A vssd1 vssd1 vccd1 vccd1 _4164_/Y sky130_fd_sc_hd__inv_2
X_4095_ _5155_/Q _4093_/C _4094_/X vssd1 vssd1 vccd1 vccd1 _4095_/Y sky130_fd_sc_hd__a21oi_1
X_3115_ _3115_/A _3115_/B vssd1 vssd1 vccd1 vccd1 _3115_/X sky130_fd_sc_hd__and2_1
X_3046_ _3106_/A _3654_/A vssd1 vssd1 vccd1 vccd1 _3046_/X sky130_fd_sc_hd__or2_1
XFILLER_36_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4997_ _5446_/CLK _4997_/D vssd1 vssd1 vccd1 vccd1 _5582_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_23_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3948_ _5263_/Q _3915_/A _3642_/B _4583_/A _3947_/X vssd1 vssd1 vccd1 vccd1 _3948_/X
+ sky130_fd_sc_hd__a221o_1
X_3879_ _3879_/A vssd1 vssd1 vccd1 vccd1 _5072_/D sky130_fd_sc_hd__clkbuf_1
X_5618_ _5618_/A _2653_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[14] sky130_fd_sc_hd__ebufn_8
X_5549_ _5549_/A _2570_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_48_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5339_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4920_ _4920_/A vssd1 vssd1 vccd1 vccd1 _5425_/D sky130_fd_sc_hd__clkbuf_1
X_4851_ _4884_/A vssd1 vssd1 vccd1 vccd1 _4851_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3802_ _5045_/Q _3803_/C _3801_/Y vssd1 vssd1 vccd1 vccd1 _5045_/D sky130_fd_sc_hd__a21oi_1
XFILLER_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4782_ _4782_/A _4782_/B vssd1 vssd1 vccd1 vccd1 _5367_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3733_ _3754_/B _3733_/B _4024_/A vssd1 vssd1 vccd1 vccd1 _3740_/A sky130_fd_sc_hd__and3_1
X_3664_ _5004_/Q _3660_/Y _3663_/X _3675_/S vssd1 vssd1 vccd1 vccd1 _5004_/D sky130_fd_sc_hd__o22a_1
X_5403_ _5445_/CLK _5403_/D vssd1 vssd1 vccd1 vccd1 _5403_/Q sky130_fd_sc_hd__dfxtp_4
X_2615_ _2616_/A vssd1 vssd1 vccd1 vccd1 _2615_/Y sky130_fd_sc_hd__inv_2
X_3595_ _5582_/A _3586_/Y _3594_/X _2761_/X vssd1 vssd1 vccd1 vccd1 _4997_/D sky130_fd_sc_hd__a211o_1
X_5334_ _5335_/CLK _5334_/D vssd1 vssd1 vccd1 vccd1 _5334_/Q sky130_fd_sc_hd__dfxtp_1
X_2546_ _2546_/A _2546_/B vssd1 vssd1 vccd1 vccd1 _5117_/D sky130_fd_sc_hd__nor2_1
X_5265_ _5323_/CLK _5265_/D vssd1 vssd1 vccd1 vccd1 _5265_/Q sky130_fd_sc_hd__dfxtp_1
X_4216_ _5418_/Q _5369_/Q _4216_/S vssd1 vssd1 vccd1 vccd1 _4216_/X sky130_fd_sc_hd__mux2_1
X_5196_ _5369_/CLK _5196_/D vssd1 vssd1 vccd1 vccd1 _5196_/Q sky130_fd_sc_hd__dfxtp_1
X_4147_ _4147_/A vssd1 vssd1 vccd1 vccd1 _5174_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4078_ _5148_/Q _2790_/B _5133_/Q vssd1 vssd1 vccd1 vccd1 _4080_/A sky130_fd_sc_hd__o21a_1
XFILLER_43_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3029_ _3029_/A _5393_/Q vssd1 vssd1 vccd1 vccd1 _3030_/B sky130_fd_sc_hd__and2_1
XFILLER_24_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3380_ _3380_/A _3380_/B vssd1 vssd1 vccd1 vccd1 _3380_/Y sky130_fd_sc_hd__nor2_1
X_5050_ _5051_/CLK _5050_/D vssd1 vssd1 vccd1 vccd1 _5050_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4903_ _5386_/D _4884_/X _4901_/Y _4902_/X vssd1 vssd1 vccd1 vccd1 _5418_/D sky130_fd_sc_hd__o211a_1
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4834_ _4834_/A _4834_/B _4834_/C _4834_/D vssd1 vssd1 vccd1 vccd1 _4835_/C sky130_fd_sc_hd__or4_1
X_4765_ _5362_/Q _5361_/Q _4765_/C vssd1 vssd1 vccd1 vccd1 _4771_/C sky130_fd_sc_hd__and3_1
X_3716_ _3750_/B vssd1 vssd1 vccd1 vccd1 _3754_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4696_ _4739_/B _4696_/B vssd1 vssd1 vccd1 vccd1 _5326_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _3647_/A _5402_/Q vssd1 vssd1 vccd1 vccd1 _3648_/B sky130_fd_sc_hd__and2_1
X_3578_ _4073_/C _3578_/B _3578_/C vssd1 vssd1 vccd1 vccd1 _3581_/B sky130_fd_sc_hd__and3_1
X_5317_ _5437_/CLK _5317_/D vssd1 vssd1 vccd1 vccd1 _5317_/Q sky130_fd_sc_hd__dfxtp_1
X_2529_ _2529_/A vssd1 vssd1 vccd1 vccd1 _5120_/D sky130_fd_sc_hd__clkbuf_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5248_ _5446_/CLK _5248_/D vssd1 vssd1 vccd1 vccd1 _5248_/Q sky130_fd_sc_hd__dfxtp_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _4000_/A _5179_/D vssd1 vssd1 vccd1 vccd1 _5179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2880_ _2849_/X _2852_/Y _3489_/B _3489_/A vssd1 vssd1 vccd1 vccd1 _5588_/A sky130_fd_sc_hd__a22o_4
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4550_ _4550_/A vssd1 vssd1 vccd1 vccd1 _5288_/D sky130_fd_sc_hd__clkbuf_1
X_4481_ _5261_/Q _5099_/Q _4481_/S vssd1 vssd1 vccd1 vccd1 _4482_/A sky130_fd_sc_hd__mux2_1
X_3501_ _5248_/Q vssd1 vssd1 vccd1 vccd1 _4730_/A sky130_fd_sc_hd__inv_2
X_3432_ _3416_/X _3431_/X _3277_/B _3260_/C vssd1 vssd1 vccd1 vccd1 _5595_/A sky130_fd_sc_hd__a211oi_2
X_3363_ _3336_/A _3380_/A _3357_/X _3267_/A _3362_/X vssd1 vssd1 vccd1 vccd1 _3363_/X
+ sky130_fd_sc_hd__a311o_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5436_/CLK _5102_/D vssd1 vssd1 vccd1 vccd1 _5102_/Q sky130_fd_sc_hd__dfxtp_1
X_3294_ _3295_/B _4074_/B _3294_/C vssd1 vssd1 vccd1 vccd1 _3396_/A sky130_fd_sc_hd__and3b_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5058_/CLK _5033_/D vssd1 vssd1 vccd1 vccd1 _5033_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4817_ _4833_/C _5398_/Q _4823_/S vssd1 vssd1 vccd1 vccd1 _4818_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4748_ _4752_/C _4748_/B vssd1 vssd1 vccd1 vccd1 _5356_/D sky130_fd_sc_hd__nor2_1
XFILLER_31_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4679_ _3892_/A _3627_/X _4586_/X _4589_/Y _4506_/Y vssd1 vssd1 vccd1 vccd1 _4680_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3981_ _5101_/Q _3976_/X _3980_/X _4833_/B vssd1 vssd1 vccd1 vccd1 _5101_/D sky130_fd_sc_hd__a22o_1
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2932_ _5304_/Q _2974_/A _2929_/X _2931_/X _2975_/A vssd1 vssd1 vccd1 vccd1 _2934_/B
+ sky130_fd_sc_hd__a221o_1
X_2863_ _5034_/Q _5033_/Q _2872_/S vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2794_ _2869_/A vssd1 vssd1 vccd1 vccd1 _2833_/A sky130_fd_sc_hd__clkbuf_2
X_5582_ _5582_/A _2609_/Y vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__ebufn_8
X_4602_ _4602_/A vssd1 vssd1 vccd1 vccd1 _5303_/D sky130_fd_sc_hd__clkbuf_1
X_4533_ _5280_/Q _5427_/Q _4541_/S vssd1 vssd1 vccd1 vccd1 _4534_/A sky130_fd_sc_hd__mux2_1
X_4464_ _5254_/Q _4674_/A _4464_/C vssd1 vssd1 vccd1 vccd1 _4471_/A sky130_fd_sc_hd__and3_1
X_3415_ _3415_/A vssd1 vssd1 vccd1 vccd1 _4902_/A sky130_fd_sc_hd__clkbuf_4
X_4395_ _5199_/Q _5169_/Q _4399_/S vssd1 vssd1 vccd1 vccd1 _4396_/B sky130_fd_sc_hd__mux2_1
X_3346_ _3372_/A _3372_/B _3345_/Y vssd1 vssd1 vccd1 vccd1 _3374_/B sky130_fd_sc_hd__o21ai_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _5058_/CLK _5016_/D vssd1 vssd1 vccd1 vccd1 _5016_/Q sky130_fd_sc_hd__dfxtp_1
X_3277_ _3424_/C _3277_/B vssd1 vssd1 vccd1 vccd1 _3277_/Y sky130_fd_sc_hd__nor2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5503__93 vssd1 vssd1 vccd1 vccd1 _5503__93/HI _5606_/A sky130_fd_sc_hd__conb_1
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3200_ _3823_/A _3823_/B _3445_/C _3191_/A vssd1 vssd1 vccd1 vccd1 _3229_/B sky130_fd_sc_hd__o31a_1
X_4180_ _4179_/X _5183_/Q _4180_/S vssd1 vssd1 vccd1 vccd1 _4181_/A sky130_fd_sc_hd__mux2_1
X_3131_ _3132_/A _3132_/B _3132_/C vssd1 vssd1 vccd1 vccd1 _3146_/B sky130_fd_sc_hd__o21a_1
X_3062_ _3118_/S vssd1 vssd1 vccd1 vccd1 _3649_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3964_ _5403_/Q _5330_/Q _4707_/B _4707_/C vssd1 vssd1 vccd1 vccd1 _4904_/C sky130_fd_sc_hd__or4_2
X_2915_ _2913_/A _2913_/B _2994_/A vssd1 vssd1 vccd1 vccd1 _2916_/B sky130_fd_sc_hd__o21ai_1
X_3895_ _3895_/A _4680_/C _4503_/B vssd1 vssd1 vccd1 vccd1 _3942_/B sky130_fd_sc_hd__nand3_1
X_5634_ _5634_/A _2673_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__ebufn_8
X_2846_ _2846_/A vssd1 vssd1 vccd1 vccd1 _2846_/X sky130_fd_sc_hd__buf_2
X_2777_ hold94/A _2717_/X _4084_/B vssd1 vssd1 vccd1 vccd1 _2778_/B sky130_fd_sc_hd__o21a_1
Xhold100 hold121/X vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__dlygate4sd3_1
X_5565_ _5565_/A _2590_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[31] sky130_fd_sc_hd__ebufn_8
Xhold122 hold89/X vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold111 hold93/X vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__clkbuf_2
Xhold144 _5095_/Q vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold133 _5084_/Q vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_4516_ _4516_/A vssd1 vssd1 vccd1 vccd1 _5272_/D sky130_fd_sc_hd__clkbuf_1
X_4447_ _4357_/A _4445_/X _4449_/B vssd1 vssd1 vccd1 vccd1 _4447_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_58_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4378_ _4667_/A vssd1 vssd1 vccd1 vccd1 _4378_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3329_ _3377_/A _3419_/B vssd1 vssd1 vccd1 vccd1 _3358_/A sky130_fd_sc_hd__and2_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2700_ _4115_/A vssd1 vssd1 vccd1 vccd1 _4708_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_9_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3680_ _4158_/A vssd1 vssd1 vccd1 vccd1 _3698_/A sky130_fd_sc_hd__buf_4
XFILLER_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2631_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2631_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5350_ _5353_/CLK _5350_/D vssd1 vssd1 vccd1 vccd1 _5350_/Q sky130_fd_sc_hd__dfxtp_1
X_2562_ _2562_/A _2562_/B vssd1 vssd1 vccd1 vccd1 _5111_/D sky130_fd_sc_hd__nor2_1
XFILLER_5_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4301_ _4300_/X _5216_/Q _4309_/S vssd1 vssd1 vccd1 vccd1 _4302_/A sky130_fd_sc_hd__mux2_1
X_5281_ _5431_/CLK _5281_/D vssd1 vssd1 vccd1 vccd1 _5281_/Q sky130_fd_sc_hd__dfxtp_1
X_4232_ _4235_/A _4232_/B vssd1 vssd1 vccd1 vccd1 _4233_/A sky130_fd_sc_hd__and2_1
XFILLER_4_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4163_ _5178_/Q _4163_/B vssd1 vssd1 vccd1 vccd1 _4164_/A sky130_fd_sc_hd__or2_1
XFILLER_55_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3114_ _3114_/A _3114_/B vssd1 vssd1 vccd1 vccd1 _3144_/B sky130_fd_sc_hd__xnor2_1
X_4094_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4094_/X sky130_fd_sc_hd__buf_4
X_5494__84 vssd1 vssd1 vccd1 vccd1 _5494__84/HI _5572_/A sky130_fd_sc_hd__conb_1
X_3045_ _3154_/A vssd1 vssd1 vccd1 vccd1 _3654_/A sky130_fd_sc_hd__buf_2
XFILLER_48_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4996_ _5439_/CLK _4996_/D vssd1 vssd1 vccd1 vccd1 _4996_/Q sky130_fd_sc_hd__dfxtp_1
X_3947_ _3947_/A vssd1 vssd1 vccd1 vccd1 _3947_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3878_ hold7/A _4834_/B _3884_/S vssd1 vssd1 vccd1 vccd1 _3879_/A sky130_fd_sc_hd__mux2_1
X_2829_ _2872_/S vssd1 vssd1 vccd1 vccd1 _2859_/S sky130_fd_sc_hd__clkbuf_2
X_5617_ _5617_/A _2652_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[13] sky130_fd_sc_hd__ebufn_8
X_5548_ _5548_/A _2569_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[14] sky130_fd_sc_hd__ebufn_8
XFILLER_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4850_ _5404_/Q _5405_/Q _5406_/Q vssd1 vssd1 vccd1 vccd1 _4855_/B sky130_fd_sc_hd__and3_1
X_3801_ _5045_/Q _3803_/C _3800_/X vssd1 vssd1 vccd1 vccd1 _3801_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_33_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4781_ _5367_/Q _4783_/C _4742_/X vssd1 vssd1 vccd1 vccd1 _4782_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3732_ _5021_/Q _3767_/A _3729_/X _3731_/Y vssd1 vssd1 vccd1 vccd1 _5021_/D sky130_fd_sc_hd__a211o_1
X_3663_ _3661_/Y _5005_/Q _5006_/Q _3662_/X _3532_/A vssd1 vssd1 vccd1 vccd1 _3663_/X
+ sky130_fd_sc_hd__o32a_1
X_5402_ _5403_/Q _5402_/D vssd1 vssd1 vccd1 vccd1 _5402_/Q sky130_fd_sc_hd__dfxtp_1
X_2614_ _2616_/A vssd1 vssd1 vccd1 vccd1 _2614_/Y sky130_fd_sc_hd__inv_2
X_3594_ _3589_/X _3593_/X _3586_/Y vssd1 vssd1 vccd1 vccd1 _3594_/X sky130_fd_sc_hd__o21ba_1
X_5333_ _5335_/CLK _5333_/D vssd1 vssd1 vccd1 vccd1 _5333_/Q sky130_fd_sc_hd__dfxtp_1
X_2545_ _5117_/Q _2541_/B _2544_/X vssd1 vssd1 vccd1 vccd1 _2546_/B sky130_fd_sc_hd__o21ai_1
X_5264_ _5437_/CLK _5264_/D vssd1 vssd1 vccd1 vccd1 _5264_/Q sky130_fd_sc_hd__dfxtp_1
X_4215_ _4215_/A vssd1 vssd1 vccd1 vccd1 _5193_/D sky130_fd_sc_hd__clkbuf_1
X_5195_ _5369_/CLK _5195_/D vssd1 vssd1 vccd1 vccd1 _5195_/Q sky130_fd_sc_hd__dfxtp_1
X_4146_ _5351_/Q _5174_/Q _4148_/S vssd1 vssd1 vccd1 vccd1 _4147_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4077_ _2760_/A _2744_/X _2750_/X vssd1 vssd1 vccd1 vccd1 _5150_/D sky130_fd_sc_hd__o21a_1
X_3028_ _3028_/A vssd1 vssd1 vccd1 vccd1 _3028_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4979_ _5452_/Q _4980_/B _4978_/X _4861_/A vssd1 vssd1 vccd1 vccd1 _5452_/D sky130_fd_sc_hd__o211a_1
XFILLER_137_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4000_ _4000_/A vssd1 vssd1 vccd1 vccd1 _4000_/X sky130_fd_sc_hd__buf_1
X_5464__54 vssd1 vssd1 vccd1 vccd1 _5464__54/HI _5541_/A sky130_fd_sc_hd__conb_1
XFILLER_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4902_ _4902_/A vssd1 vssd1 vccd1 vccd1 _4902_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4833_ _4833_/A _4833_/B _4833_/C _4833_/D vssd1 vssd1 vccd1 vccd1 _4834_/D sky130_fd_sc_hd__or4_1
X_4764_ _4764_/A _4764_/B vssd1 vssd1 vccd1 vccd1 _5361_/D sky130_fd_sc_hd__nor2_1
X_3715_ _3715_/A vssd1 vssd1 vccd1 vccd1 _3734_/B sky130_fd_sc_hd__clkbuf_2
X_4695_ _4698_/B _4693_/Y _4694_/Y _4588_/X _4586_/C vssd1 vssd1 vccd1 vccd1 _4696_/B
+ sky130_fd_sc_hd__o32a_1
X_3646_ _3646_/A _3646_/B _3646_/C vssd1 vssd1 vccd1 vccd1 _3655_/A sky130_fd_sc_hd__or3_2
XFILLER_136_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3577_ _3577_/A _3577_/B vssd1 vssd1 vccd1 vccd1 _4993_/D sky130_fd_sc_hd__nor2_1
X_5316_ _5437_/CLK _5316_/D vssd1 vssd1 vccd1 vccd1 _5316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2528_ _2530_/B _2560_/B vssd1 vssd1 vccd1 vccd1 _2529_/A sky130_fd_sc_hd__and2_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5247_ _4000_/A _5247_/D vssd1 vssd1 vccd1 vccd1 _5247_/Q sky130_fd_sc_hd__dfxtp_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _5245_/CLK _5178_/D vssd1 vssd1 vccd1 vccd1 _5178_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4129_ _5343_/Q _5166_/Q _4137_/S vssd1 vssd1 vccd1 vccd1 _4130_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3500_ _3662_/C vssd1 vssd1 vccd1 vccd1 _4432_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4480_ _4480_/A vssd1 vssd1 vccd1 vccd1 _5260_/D sky130_fd_sc_hd__clkbuf_1
X_3431_ _3431_/A _4075_/B _3430_/X vssd1 vssd1 vccd1 vccd1 _3431_/X sky130_fd_sc_hd__or3b_1
X_3362_ _3418_/S _3344_/X _3343_/A vssd1 vssd1 vccd1 vccd1 _3362_/X sky130_fd_sc_hd__o21a_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5436_/CLK _5101_/D vssd1 vssd1 vccd1 vccd1 _5101_/Q sky130_fd_sc_hd__dfxtp_1
X_3293_ _4994_/Q _3438_/B vssd1 vssd1 vccd1 vccd1 _3294_/C sky130_fd_sc_hd__or2_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5032_/CLK _5032_/D vssd1 vssd1 vccd1 vccd1 _5032_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_10_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5313_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_26_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4816_ _4816_/A vssd1 vssd1 vccd1 vccd1 _5397_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4747_ _5356_/Q _4744_/A _4746_/X vssd1 vssd1 vccd1 vccd1 _4748_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4678_ _4594_/A _4681_/A _3945_/B _4508_/B vssd1 vssd1 vccd1 vccd1 _4678_/X sky130_fd_sc_hd__a31o_1
X_3629_ _5002_/Q vssd1 vssd1 vccd1 vccd1 _3642_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ _3980_/A vssd1 vssd1 vccd1 vccd1 _3980_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _5601_/A _4964_/A _2930_/X _2953_/C vssd1 vssd1 vccd1 vccd1 _2931_/X sky130_fd_sc_hd__a22o_1
XFILLER_30_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2862_ _2857_/X _2860_/X _4034_/A vssd1 vssd1 vccd1 vccd1 _2862_/X sky130_fd_sc_hd__mux2_1
X_4601_ _4609_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4602_/A sky130_fd_sc_hd__and2_1
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2793_ _5127_/Q vssd1 vssd1 vccd1 vccd1 _2869_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5581_ _5581_/A _2608_/Y vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__ebufn_8
XFILLER_30_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4532_ _4532_/A vssd1 vssd1 vccd1 vccd1 _4541_/S sky130_fd_sc_hd__clkbuf_2
X_4463_ _4504_/A _4504_/B vssd1 vssd1 vccd1 vccd1 _4464_/C sky130_fd_sc_hd__and2b_1
X_3414_ _3396_/Y _3399_/Y _3409_/X _3413_/Y _3305_/B vssd1 vssd1 vccd1 vccd1 _3414_/X
+ sky130_fd_sc_hd__o2111a_1
X_4394_ _3649_/A _4383_/X _4393_/X _4378_/X vssd1 vssd1 vccd1 vccd1 _5235_/D sky130_fd_sc_hd__o211a_1
X_3345_ _3337_/B _3344_/X _3337_/A vssd1 vssd1 vccd1 vccd1 _3345_/Y sky130_fd_sc_hd__a21oi_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _5056_/Q vssd1 vssd1 vccd1 vccd1 _3424_/C sky130_fd_sc_hd__clkbuf_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5058_/CLK _5015_/D vssd1 vssd1 vccd1 vccd1 _5015_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3130_ _3130_/A _3130_/B vssd1 vssd1 vccd1 vccd1 _3132_/C sky130_fd_sc_hd__xnor2_1
XFILLER_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3061_ _3084_/A vssd1 vssd1 vccd1 vccd1 _3118_/S sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3963_ _5333_/Q _5335_/Q _5334_/Q vssd1 vssd1 vccd1 vccd1 _4707_/C sky130_fd_sc_hd__or3b_1
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_3894_ _3912_/A _3894_/B vssd1 vssd1 vccd1 vccd1 _4503_/B sky130_fd_sc_hd__nand2_1
X_2914_ _5235_/Q vssd1 vssd1 vccd1 vccd1 _2994_/A sky130_fd_sc_hd__clkbuf_2
X_5633_ _5633_/A _2671_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__ebufn_8
X_2845_ _2860_/S vssd1 vssd1 vccd1 vccd1 _2846_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_12_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5564_ _5564_/A _2589_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[30] sky130_fd_sc_hd__ebufn_8
Xhold101 hold120/X vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__clkbuf_2
X_2776_ _5151_/Q vssd1 vssd1 vccd1 vccd1 _4084_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4515_ _4515_/A _4515_/B _4515_/C vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__or3_1
Xhold123 hold88/X vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold112 hold92/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__clkbuf_1
Xhold134 _5182_/Q vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_4446_ _4449_/B _4357_/A _3682_/B _3529_/A vssd1 vssd1 vccd1 vccd1 _4446_/X sky130_fd_sc_hd__a22o_1
X_4377_ _4634_/A vssd1 vssd1 vccd1 vccd1 _4667_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3328_ _3328_/A vssd1 vssd1 vccd1 vccd1 _3419_/B sky130_fd_sc_hd__clkbuf_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _3572_/B _3260_/D _3396_/B vssd1 vssd1 vccd1 vccd1 _3305_/B sky130_fd_sc_hd__o21bai_2
XFILLER_27_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2630_ _2634_/A vssd1 vssd1 vccd1 vccd1 _2630_/Y sky130_fd_sc_hd__inv_2
X_2561_ _3705_/B _2564_/A _2544_/X vssd1 vssd1 vccd1 vccd1 _2562_/B sky130_fd_sc_hd__o21ai_1
XFILLER_5_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4300_ _5212_/Q _4264_/X _4299_/X vssd1 vssd1 vccd1 vccd1 _4300_/X sky130_fd_sc_hd__a21o_1
X_5280_ _5430_/CLK _5280_/D vssd1 vssd1 vccd1 vccd1 _5280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4231_ _5198_/Q input9/X _4234_/S vssd1 vssd1 vccd1 vccd1 _4232_/B sky130_fd_sc_hd__mux2_1
X_4162_ _4112_/A _4163_/B _4161_/Y vssd1 vssd1 vccd1 vccd1 _5177_/D sky130_fd_sc_hd__o21ai_1
X_4093_ _4093_/A _4093_/B _4093_/C vssd1 vssd1 vccd1 vccd1 _5154_/D sky130_fd_sc_hd__nor3_1
X_3113_ _3114_/A _3114_/B vssd1 vssd1 vccd1 vccd1 _3146_/A sky130_fd_sc_hd__or2_1
XFILLER_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3044_ _3134_/A vssd1 vssd1 vccd1 vccd1 _3154_/A sky130_fd_sc_hd__buf_6
XFILLER_24_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4995_ _5439_/CLK _4995_/D vssd1 vssd1 vccd1 vccd1 _4995_/Q sky130_fd_sc_hd__dfxtp_1
X_5530__120 vssd1 vssd1 vccd1 vccd1 _5530__120/HI _5530__120/LO sky130_fd_sc_hd__conb_1
XFILLER_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3946_ _3946_/A _3946_/B vssd1 vssd1 vccd1 vccd1 _3947_/A sky130_fd_sc_hd__and2_1
XFILLER_32_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3877_ _3877_/A vssd1 vssd1 vccd1 vccd1 _5071_/D sky130_fd_sc_hd__clkbuf_1
X_2828_ _3474_/B vssd1 vssd1 vccd1 vccd1 _3480_/B sky130_fd_sc_hd__clkbuf_2
X_5616_ _5617_/A _2651_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[12] sky130_fd_sc_hd__ebufn_8
X_5547_ _5547_/A _2568_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[13] sky130_fd_sc_hd__ebufn_8
X_2759_ _2759_/A _5040_/Q vssd1 vssd1 vccd1 vccd1 _2759_/X sky130_fd_sc_hd__or2b_1
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4429_ _4165_/A _4115_/B _4436_/A vssd1 vssd1 vccd1 vccd1 _4429_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_48_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5514__104 vssd1 vssd1 vccd1 vccd1 _5514__104/HI _5625_/A sky130_fd_sc_hd__conb_1
XFILLER_33_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4780_ _5367_/Q _5366_/Q _4780_/C vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__and3_1
X_3800_ _3805_/C vssd1 vssd1 vccd1 vccd1 _3800_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3731_ _3720_/B _3730_/X _3729_/B vssd1 vssd1 vccd1 vccd1 _3731_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_13_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3662_ _5248_/Q _3673_/B _3662_/C vssd1 vssd1 vccd1 vccd1 _3662_/X sky130_fd_sc_hd__and3_1
X_5401_ _5403_/Q _5401_/D vssd1 vssd1 vccd1 vccd1 _5401_/Q sky130_fd_sc_hd__dfxtp_1
X_3593_ _5219_/Q _3534_/B _3541_/X _5173_/Q _3592_/Y vssd1 vssd1 vccd1 vccd1 _3593_/X
+ sky130_fd_sc_hd__a221o_1
X_2613_ _2616_/A vssd1 vssd1 vccd1 vccd1 _2613_/Y sky130_fd_sc_hd__inv_2
X_2544_ _2548_/C vssd1 vssd1 vccd1 vccd1 _2544_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5332_ _5335_/CLK _5332_/D vssd1 vssd1 vccd1 vccd1 _5332_/Q sky130_fd_sc_hd__dfxtp_1
X_5263_ _5435_/CLK _5263_/D vssd1 vssd1 vccd1 vccd1 _5263_/Q sky130_fd_sc_hd__dfxtp_1
X_5194_ _5351_/CLK _5194_/D vssd1 vssd1 vccd1 vccd1 _5194_/Q sky130_fd_sc_hd__dfxtp_1
X_4214_ _4213_/X _5193_/Q _4214_/S vssd1 vssd1 vccd1 vccd1 _4215_/A sky130_fd_sc_hd__mux2_1
X_4145_ _4145_/A vssd1 vssd1 vccd1 vccd1 _5173_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3998__6 _3999__7/A vssd1 vssd1 vccd1 vccd1 _5113_/CLK sky130_fd_sc_hd__inv_2
XFILLER_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4076_ hold135/X _4024_/A _4075_/X vssd1 vssd1 vccd1 vccd1 _5149_/D sky130_fd_sc_hd__a21bo_1
X_3027_ _3027_/A vssd1 vssd1 vccd1 vccd1 _3028_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4978_ _4978_/A _4982_/B vssd1 vssd1 vccd1 vccd1 _4978_/X sky130_fd_sc_hd__or2_1
X_3929_ _5259_/Q _3919_/X _3897_/X _5081_/Q vssd1 vssd1 vccd1 vccd1 _3929_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4901_ _4901_/A _4901_/B vssd1 vssd1 vccd1 vccd1 _4901_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4832_ _4832_/A _4832_/B _4832_/C _4832_/D vssd1 vssd1 vccd1 vccd1 _4833_/D sky130_fd_sc_hd__or4_1
XFILLER_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4763_ _5361_/Q _4765_/C _4762_/X vssd1 vssd1 vccd1 vccd1 _4764_/B sky130_fd_sc_hd__o21ai_1
X_3714_ _3710_/X _3713_/X _5016_/Q _3711_/X vssd1 vssd1 vccd1 vccd1 _5016_/D sky130_fd_sc_hd__o2bb2a_1
X_4694_ _5326_/Q _4694_/B vssd1 vssd1 vccd1 vccd1 _4694_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3645_ _5003_/Q vssd1 vssd1 vccd1 vccd1 _3645_/Y sky130_fd_sc_hd__inv_2
XFILLER_136_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3576_ _3551_/C _3574_/A _3569_/X vssd1 vssd1 vccd1 vccd1 _3577_/B sky130_fd_sc_hd__o21ai_1
X_5315_ _5328_/CLK _5315_/D vssd1 vssd1 vccd1 vccd1 _5315_/Q sky130_fd_sc_hd__dfxtp_1
X_2527_ _5587_/A _2527_/B vssd1 vssd1 vccd1 vccd1 _2560_/B sky130_fd_sc_hd__nor2_1
X_5246_ _5446_/CLK _5246_/D vssd1 vssd1 vccd1 vccd1 _5246_/Q sky130_fd_sc_hd__dfxtp_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _5245_/CLK _5177_/D vssd1 vssd1 vccd1 vccd1 _5177_/Q sky130_fd_sc_hd__dfxtp_1
X_4128_ _4261_/S vssd1 vssd1 vccd1 vccd1 _4137_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4059_ _5378_/Q hold52/A _4065_/S vssd1 vssd1 vccd1 vccd1 _4060_/A sky130_fd_sc_hd__mux2_1
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3430_ _4074_/B _3396_/B _3429_/X _3415_/A vssd1 vssd1 vccd1 vccd1 _3430_/X sky130_fd_sc_hd__o211a_1
X_3361_ _3343_/A _3359_/X _3390_/A _3360_/Y vssd1 vssd1 vccd1 vccd1 _3361_/X sky130_fd_sc_hd__a31o_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5436_/CLK _5100_/D vssd1 vssd1 vccd1 vccd1 _5100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5031_ _5032_/CLK _5031_/D vssd1 vssd1 vccd1 vccd1 _5031_/Q sky130_fd_sc_hd__dfxtp_1
X_3292_ _3292_/A vssd1 vssd1 vccd1 vccd1 _4074_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_2_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4815_ _4834_/B _5397_/Q _4823_/S vssd1 vssd1 vccd1 vccd1 _4816_/A sky130_fd_sc_hd__mux2_1
X_4746_ _4762_/A vssd1 vssd1 vccd1 vccd1 _4746_/X sky130_fd_sc_hd__clkbuf_2
X_4677_ _5320_/Q _4676_/X _4583_/B _4093_/A vssd1 vssd1 vccd1 vccd1 _5320_/D sky130_fd_sc_hd__a211o_1
X_3628_ _5323_/Q _4328_/A _5321_/Q vssd1 vssd1 vccd1 vccd1 _3892_/B sky130_fd_sc_hd__or3_2
X_3559_ _4789_/B _3559_/B _3559_/C vssd1 vssd1 vccd1 vccd1 _3560_/A sky130_fd_sc_hd__and3_1
X_5229_ _5445_/CLK _5229_/D vssd1 vssd1 vccd1 vccd1 _5229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_48_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2930_ _5452_/Q _5372_/Q vssd1 vssd1 vccd1 vccd1 _2930_/X sky130_fd_sc_hd__or2b_1
XFILLER_15_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2861_ _3464_/A vssd1 vssd1 vccd1 vccd1 _4034_/A sky130_fd_sc_hd__clkbuf_2
X_4600_ _5303_/Q _4596_/X _4617_/S vssd1 vssd1 vccd1 vccd1 _4601_/B sky130_fd_sc_hd__mux2_1
X_2792_ _3888_/S vssd1 vssd1 vccd1 vccd1 _5133_/D sky130_fd_sc_hd__buf_2
X_5580_ _5580_/A _2607_/Y vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__ebufn_8
X_4531_ _4531_/A vssd1 vssd1 vccd1 vccd1 _5279_/D sky130_fd_sc_hd__clkbuf_1
X_4462_ _5436_/Q _5437_/Q _3415_/A vssd1 vssd1 vccd1 vccd1 _4674_/A sky130_fd_sc_hd__o21a_1
X_3413_ _3413_/A _3413_/B vssd1 vssd1 vccd1 vccd1 _3413_/Y sky130_fd_sc_hd__xnor2_1
X_4393_ _4400_/A _4393_/B vssd1 vssd1 vccd1 vccd1 _4393_/X sky130_fd_sc_hd__or2_1
X_3344_ _3344_/A vssd1 vssd1 vccd1 vccd1 _3344_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3275_/A _3275_/B vssd1 vssd1 vccd1 vccd1 _3280_/B sky130_fd_sc_hd__nor2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5014_ _5431_/CLK _5014_/D vssd1 vssd1 vccd1 vccd1 _5014_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4729_ hold139/X _4727_/A _4728_/Y vssd1 vssd1 vccd1 vccd1 _5335_/D sky130_fd_sc_hd__a21oi_1
XFILLER_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3060_ _3060_/A _3060_/B vssd1 vssd1 vccd1 vccd1 _4832_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3962_ _5329_/Q _5332_/Q _5331_/Q vssd1 vssd1 vccd1 vccd1 _4707_/B sky130_fd_sc_hd__or3_1
X_2913_ _2913_/A _2913_/B vssd1 vssd1 vccd1 vccd1 _2939_/A sky130_fd_sc_hd__nand2_1
X_3893_ _4504_/A _3893_/B vssd1 vssd1 vccd1 vccd1 _3894_/B sky130_fd_sc_hd__nor2_1
X_5632_ _5632_/A _2670_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__ebufn_8
X_2844_ _5033_/Q _3480_/B vssd1 vssd1 vccd1 vccd1 _2844_/X sky130_fd_sc_hd__and2_1
X_5563_ _5563_/A _2588_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[29] sky130_fd_sc_hd__ebufn_8
X_2775_ _2889_/B _4959_/B _3967_/A _2889_/A vssd1 vssd1 vccd1 vccd1 _2775_/X sky130_fd_sc_hd__or4b_2
X_4514_ _4551_/B _4514_/B vssd1 vssd1 vccd1 vccd1 _4515_/C sky130_fd_sc_hd__nor2_1
Xhold124 hold95/X vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold113 _5155_/Q vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold102 _5064_/Q vssd1 vssd1 vccd1 vccd1 hold129/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _5149_/Q vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_4445_ _4450_/B vssd1 vssd1 vccd1 vccd1 _4445_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4376_ _4381_/A _4376_/B vssd1 vssd1 vccd1 vccd1 _4376_/X sky130_fd_sc_hd__or2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _4987_/Q vssd1 vssd1 vccd1 vccd1 _3377_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _3438_/B _3398_/A _3260_/C vssd1 vssd1 vccd1 vccd1 _3396_/B sky130_fd_sc_hd__a21oi_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3189_ _5053_/Q vssd1 vssd1 vccd1 vccd1 _3445_/C sky130_fd_sc_hd__inv_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2560_ _3705_/C _2560_/B vssd1 vssd1 vccd1 vccd1 _2564_/A sky130_fd_sc_hd__and2_1
X_4230_ _4230_/A vssd1 vssd1 vccd1 vccd1 _5197_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_4_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4161_ _4161_/A _4161_/B vssd1 vssd1 vccd1 vccd1 _4161_/Y sky130_fd_sc_hd__nand2_1
X_4092_ _4092_/A _4092_/B vssd1 vssd1 vccd1 vccd1 _4093_/C sky130_fd_sc_hd__and2_1
X_3112_ _3142_/A _3112_/B vssd1 vssd1 vccd1 vccd1 _3114_/B sky130_fd_sc_hd__xnor2_1
X_3043_ _3134_/A _3043_/B vssd1 vssd1 vccd1 vccd1 _4833_/A sky130_fd_sc_hd__xnor2_4
XFILLER_36_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4994_ _5335_/CLK _4994_/D vssd1 vssd1 vccd1 vccd1 _4994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3945_ _5324_/Q _3945_/B vssd1 vssd1 vccd1 vccd1 _3946_/B sky130_fd_sc_hd__nand2_1
X_3876_ hold1/A _4834_/A _3884_/S vssd1 vssd1 vccd1 vccd1 _3877_/A sky130_fd_sc_hd__mux2_1
X_5615_ _5617_/A _2650_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[11] sky130_fd_sc_hd__ebufn_8
X_2827_ _2840_/A _5132_/Q _2827_/C vssd1 vssd1 vccd1 vccd1 _3474_/B sky130_fd_sc_hd__or3_1
X_5546_ _5546_/A _2682_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[12] sky130_fd_sc_hd__ebufn_8
X_2758_ _2753_/Y _2755_/X _4739_/B vssd1 vssd1 vccd1 vccd1 _5039_/D sky130_fd_sc_hd__a21oi_1
X_2689_ _2689_/A vssd1 vssd1 vccd1 vccd1 _2689_/Y sky130_fd_sc_hd__inv_2
X_4428_ _4428_/A vssd1 vssd1 vccd1 vccd1 _5244_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4359_ _5227_/Q _4350_/X _4353_/X _5249_/D vssd1 vssd1 vccd1 vccd1 _5227_/D sky130_fd_sc_hd__a22o_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5058_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5485__75 vssd1 vssd1 vccd1 vccd1 _5485__75/HI _5563_/A sky130_fd_sc_hd__conb_1
XFILLER_27_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3730_ _3709_/B _3754_/B _3750_/A vssd1 vssd1 vccd1 vccd1 _3730_/X sky130_fd_sc_hd__a21bo_1
XFILLER_13_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3661_ _5004_/Q vssd1 vssd1 vccd1 vccd1 _3661_/Y sky130_fd_sc_hd__inv_2
X_5400_ _5403_/Q _5400_/D vssd1 vssd1 vccd1 vccd1 _5400_/Q sky130_fd_sc_hd__dfxtp_1
X_3592_ _3592_/A _4434_/B _3592_/C vssd1 vssd1 vccd1 vccd1 _3592_/Y sky130_fd_sc_hd__nor3_1
X_2612_ _2616_/A vssd1 vssd1 vccd1 vccd1 _2612_/Y sky130_fd_sc_hd__inv_2
X_2543_ _3705_/A _2546_/A _2542_/Y vssd1 vssd1 vccd1 vccd1 _5118_/D sky130_fd_sc_hd__o21a_1
X_5331_ _5446_/CLK _5331_/D vssd1 vssd1 vccd1 vccd1 _5331_/Q sky130_fd_sc_hd__dfxtp_1
X_5262_ _5435_/CLK _5262_/D vssd1 vssd1 vccd1 vccd1 _5262_/Q sky130_fd_sc_hd__dfxtp_1
X_5193_ _5369_/CLK _5193_/D vssd1 vssd1 vccd1 vccd1 _5193_/Q sky130_fd_sc_hd__dfxtp_1
X_4213_ _5417_/Q _5368_/Q _4216_/S vssd1 vssd1 vccd1 vccd1 _4213_/X sky130_fd_sc_hd__mux2_1
X_4144_ _5350_/Q _5173_/Q _4148_/S vssd1 vssd1 vccd1 vccd1 _4145_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4075_ _4075_/A _4075_/B _4075_/C _4075_/D vssd1 vssd1 vccd1 vccd1 _4075_/X sky130_fd_sc_hd__or4_1
X_3026_ _2944_/X _4832_/B _3025_/X vssd1 vssd1 vccd1 vccd1 _5377_/D sky130_fd_sc_hd__o21a_1
XFILLER_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4977_ input15/X _4982_/B _4976_/X _4861_/A vssd1 vssd1 vccd1 vccd1 _5451_/D sky130_fd_sc_hd__o211a_1
XFILLER_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3928_ hold143/X _3909_/X _3927_/X vssd1 vssd1 vccd1 vccd1 _5084_/D sky130_fd_sc_hd__o21a_1
XFILLER_137_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3859_ _3859_/A vssd1 vssd1 vccd1 vccd1 _5063_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ _5418_/Q _4900_/B vssd1 vssd1 vccd1 vccd1 _4901_/B sky130_fd_sc_hd__xor2_1
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4831_ _4831_/A _4831_/B _4831_/C _4831_/D vssd1 vssd1 vccd1 vccd1 _4832_/D sky130_fd_sc_hd__or4_1
X_4762_ _4762_/A vssd1 vssd1 vccd1 vccd1 _4762_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3713_ _3726_/A _3726_/B _3713_/C_N vssd1 vssd1 vccd1 vccd1 _3713_/X sky130_fd_sc_hd__or3b_1
X_4693_ _4693_/A _4693_/B vssd1 vssd1 vccd1 vccd1 _4693_/Y sky130_fd_sc_hd__nand2_1
X_3644_ _3644_/A vssd1 vssd1 vccd1 vccd1 _5002_/D sky130_fd_sc_hd__clkbuf_1
X_3575_ _3578_/B _3575_/B vssd1 vssd1 vccd1 vccd1 _3577_/A sky130_fd_sc_hd__and2_1
X_5314_ _5328_/CLK _5314_/D vssd1 vssd1 vccd1 vccd1 _5314_/Q sky130_fd_sc_hd__dfxtp_1
X_2526_ _2548_/C vssd1 vssd1 vccd1 vccd1 _2530_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5245_ _5245_/CLK _5245_/D vssd1 vssd1 vccd1 vccd1 _5245_/Q sky130_fd_sc_hd__dfxtp_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5176_ _5339_/CLK _5176_/D vssd1 vssd1 vccd1 vccd1 _5176_/Q sky130_fd_sc_hd__dfxtp_1
X_4127_ _4127_/A vssd1 vssd1 vccd1 vccd1 _5165_/D sky130_fd_sc_hd__clkbuf_1
X_4058_ _4058_/A vssd1 vssd1 vccd1 vccd1 _5140_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5456__125 vssd1 vssd1 vccd1 vccd1 _5456__125/HI _5456__125/LO sky130_fd_sc_hd__conb_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3009_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3009_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3360_ _3563_/A _3551_/B _3334_/A _3267_/A vssd1 vssd1 vccd1 vccd1 _3360_/Y sky130_fd_sc_hd__o31ai_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5032_/CLK _5030_/D vssd1 vssd1 vccd1 vccd1 _5030_/Q sky130_fd_sc_hd__dfxtp_1
X_3291_ _3318_/A _3313_/B vssd1 vssd1 vccd1 vccd1 _3411_/A sky130_fd_sc_hd__and2b_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4814_ _4825_/S vssd1 vssd1 vccd1 vccd1 _4823_/S sky130_fd_sc_hd__clkbuf_2
X_4745_ _5356_/Q _5355_/Q _5371_/D vssd1 vssd1 vccd1 vccd1 _4752_/C sky130_fd_sc_hd__and3_1
XFILLER_21_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4676_ _5301_/Q _3915_/X _4508_/B _4675_/Y vssd1 vssd1 vccd1 vccd1 _4676_/X sky130_fd_sc_hd__a211o_1
X_3627_ _3895_/A vssd1 vssd1 vccd1 vccd1 _3627_/X sky130_fd_sc_hd__buf_2
X_3558_ _3563_/C vssd1 vssd1 vccd1 vccd1 _3559_/C sky130_fd_sc_hd__clkinv_2
XFILLER_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3489_ _3489_/A _3489_/B vssd1 vssd1 vccd1 vccd1 _3490_/A sky130_fd_sc_hd__or2_4
X_5228_ _5445_/CLK _5228_/D vssd1 vssd1 vccd1 vccd1 _5228_/Q sky130_fd_sc_hd__dfxtp_1
X_5159_ _5160_/CLK _5159_/D vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2860_ _2858_/X _2859_/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2860_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2791_ _4044_/A vssd1 vssd1 vccd1 vccd1 _3888_/S sky130_fd_sc_hd__clkinv_2
XFILLER_31_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4530_ _5279_/Q _5426_/Q _4530_/S vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__mux2_1
XFILLER_7_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4461_ _4739_/B _4693_/A vssd1 vssd1 vccd1 vccd1 _5254_/D sky130_fd_sc_hd__nor2_1
X_3412_ _3412_/A _3412_/B vssd1 vssd1 vccd1 vccd1 _3413_/B sky130_fd_sc_hd__nor2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4392_ _5198_/Q _5168_/Q _4399_/S vssd1 vssd1 vccd1 vccd1 _4393_/B sky130_fd_sc_hd__mux2_1
X_3343_ _3343_/A _3343_/B vssd1 vssd1 vccd1 vccd1 _3372_/B sky130_fd_sc_hd__nand2_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _3309_/A _3307_/B vssd1 vssd1 vccd1 vccd1 _3300_/A sky130_fd_sc_hd__nand2b_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5430_/CLK _5013_/D vssd1 vssd1 vccd1 vccd1 _5013_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2989_ _3023_/A _2989_/B vssd1 vssd1 vccd1 vccd1 _4831_/D sky130_fd_sc_hd__xor2_1
X_4728_ _5335_/Q _4727_/A _4710_/B vssd1 vssd1 vccd1 vccd1 _4728_/Y sky130_fd_sc_hd__o21ai_1
X_4659_ _4667_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4660_/A sky130_fd_sc_hd__and2_1
XFILLER_49_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5051_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_51_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3961_ _5419_/Q vssd1 vssd1 vccd1 vccd1 _3961_/Y sky130_fd_sc_hd__inv_2
X_2912_ _3033_/A _2912_/B vssd1 vssd1 vccd1 vccd1 _2913_/B sky130_fd_sc_hd__xnor2_2
X_3892_ _3892_/A _3892_/B vssd1 vssd1 vccd1 vccd1 _4680_/C sky130_fd_sc_hd__or2_1
X_5631_ _5631_/A _2669_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__ebufn_8
X_2843_ _2841_/X _2842_/X _2843_/S vssd1 vssd1 vccd1 vccd1 _2843_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5562_ _5562_/A _2587_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[28] sky130_fd_sc_hd__ebufn_8
X_2774_ _5386_/Q vssd1 vssd1 vccd1 vccd1 _2889_/A sky130_fd_sc_hd__clkbuf_4
X_4513_ _5271_/Q _4514_/B _5272_/Q vssd1 vssd1 vccd1 vccd1 _4515_/B sky130_fd_sc_hd__o21a_1
Xhold114 hold97/X vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__clkbuf_2
Xhold125 hold94/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold103 hold129/X vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__clkbuf_2
X_4444_ _4165_/A _4438_/B _4443_/Y _4350_/X vssd1 vssd1 vccd1 vccd1 _5248_/D sky130_fd_sc_hd__o211ai_1
X_4375_ input9/X _5164_/Q _4380_/S vssd1 vssd1 vccd1 vccd1 _4376_/B sky130_fd_sc_hd__mux2_1
X_3326_ _4988_/Q vssd1 vssd1 vccd1 vccd1 _4073_/D sky130_fd_sc_hd__clkbuf_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3295_/B _3292_/A vssd1 vssd1 vccd1 vccd1 _3260_/C sky130_fd_sc_hd__nor2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3188_ _2889_/A _3028_/A _3186_/X _3120_/X _3187_/X vssd1 vssd1 vccd1 vccd1 _5386_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_27_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4160_ _5177_/Q _4161_/B vssd1 vssd1 vccd1 vccd1 _4163_/B sky130_fd_sc_hd__or2_1
X_3111_ _3129_/A _3111_/B vssd1 vssd1 vccd1 vccd1 _3112_/B sky130_fd_sc_hd__and2_1
XFILLER_4_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4091_ _2781_/B _4092_/B _5154_/Q vssd1 vssd1 vccd1 vccd1 _4093_/B sky130_fd_sc_hd__a21oi_1
X_3042_ _3036_/A _3040_/Y _3084_/A vssd1 vssd1 vccd1 vccd1 _3043_/B sky130_fd_sc_hd__mux2_2
XFILLER_48_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4993_ _5446_/CLK _4993_/D vssd1 vssd1 vccd1 vccd1 _4993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3944_ _5301_/Q vssd1 vssd1 vccd1 vccd1 _4583_/A sky130_fd_sc_hd__inv_2
X_3875_ _3888_/S vssd1 vssd1 vccd1 vccd1 _3884_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_137_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2826_ _2826_/A vssd1 vssd1 vccd1 vccd1 _3466_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5614_ _5617_/A _2649_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[10] sky130_fd_sc_hd__ebufn_8
XFILLER_31_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2757_ _4685_/A vssd1 vssd1 vccd1 vccd1 _4739_/B sky130_fd_sc_hd__buf_4
X_5545_ _5545_/A _2692_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[11] sky130_fd_sc_hd__ebufn_8
X_2688_ _2689_/A vssd1 vssd1 vccd1 vccd1 _2688_/Y sky130_fd_sc_hd__inv_2
X_4427_ _4685_/A _4427_/B vssd1 vssd1 vccd1 vccd1 _4428_/A sky130_fd_sc_hd__or2_1
XFILLER_59_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _4357_/A _4356_/X _4357_/Y _4350_/A vssd1 vssd1 vccd1 vccd1 _5249_/D sky130_fd_sc_hd__o211a_1
X_3309_ _3309_/A _3309_/B vssd1 vssd1 vccd1 vccd1 _3309_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4289_ _4289_/A vssd1 vssd1 vccd1 vccd1 _5213_/D sky130_fd_sc_hd__clkbuf_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4007__2 _5439_/CLK vssd1 vssd1 vccd1 vccd1 _5121_/CLK sky130_fd_sc_hd__inv_2
XFILLER_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3660_ _5005_/Q _3675_/S vssd1 vssd1 vccd1 vccd1 _3660_/Y sky130_fd_sc_hd__nor2_1
X_3591_ _4449_/B _4449_/C _3510_/C _5251_/Q vssd1 vssd1 vccd1 vccd1 _3592_/C sky130_fd_sc_hd__o211a_1
X_2611_ _2635_/A vssd1 vssd1 vccd1 vccd1 _2616_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2542_ _3705_/A _2546_/A _2530_/B vssd1 vssd1 vccd1 vccd1 _2542_/Y sky130_fd_sc_hd__a21boi_1
X_5330_ _5446_/CLK _5330_/D vssd1 vssd1 vccd1 vccd1 _5330_/Q sky130_fd_sc_hd__dfxtp_1
X_5261_ _5435_/CLK _5261_/D vssd1 vssd1 vccd1 vccd1 _5261_/Q sky130_fd_sc_hd__dfxtp_1
X_4212_ _4212_/A vssd1 vssd1 vccd1 vccd1 _5192_/D sky130_fd_sc_hd__clkbuf_1
X_5192_ _5369_/CLK _5192_/D vssd1 vssd1 vccd1 vccd1 _5192_/Q sky130_fd_sc_hd__dfxtp_1
X_4143_ _4143_/A vssd1 vssd1 vccd1 vccd1 _5172_/D sky130_fd_sc_hd__clkbuf_1
X_4074_ _4115_/A _4074_/B _4073_/X _2760_/A vssd1 vssd1 vccd1 vccd1 _4075_/D sky130_fd_sc_hd__or4bb_1
X_3025_ _2991_/A _5377_/Q _5233_/Q vssd1 vssd1 vccd1 vccd1 _3025_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4976_ _5451_/Q _4980_/B vssd1 vssd1 vccd1 vccd1 _4976_/X sky130_fd_sc_hd__or2_1
X_3927_ _5284_/Q _3910_/X _3697_/A _3926_/X vssd1 vssd1 vccd1 vccd1 _3927_/X sky130_fd_sc_hd__a211o_1
XFILLER_137_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3858_ _5063_/Q _2942_/X _5133_/D vssd1 vssd1 vccd1 vccd1 _3859_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2809_ _5127_/Q vssd1 vssd1 vccd1 vccd1 _2872_/S sky130_fd_sc_hd__clkbuf_2
X_3789_ _3789_/A vssd1 vssd1 vccd1 vccd1 _5041_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5520__110 vssd1 vssd1 vccd1 vccd1 _5520__110/HI _5636_/A sky130_fd_sc_hd__conb_1
XFILLER_49_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4830_ _4830_/A vssd1 vssd1 vccd1 vccd1 _5403_/D sky130_fd_sc_hd__clkbuf_1
X_4761_ _5361_/Q _4765_/C vssd1 vssd1 vccd1 vccd1 _4764_/A sky130_fd_sc_hd__and2_1
X_3712_ _3707_/X _3710_/X _5015_/Q _3711_/X vssd1 vssd1 vccd1 vccd1 _5015_/D sky130_fd_sc_hd__o2bb2a_1
X_4692_ _5326_/Q _4692_/B _4692_/C vssd1 vssd1 vccd1 vccd1 _4698_/B sky130_fd_sc_hd__and3_1
X_3643_ _3642_/Y _3642_/A _3643_/S vssd1 vssd1 vccd1 vccd1 _3644_/A sky130_fd_sc_hd__mux2_1
X_5313_ _5313_/CLK _5313_/D vssd1 vssd1 vccd1 vccd1 _5313_/Q sky130_fd_sc_hd__dfxtp_1
X_3574_ _3574_/A _3574_/B vssd1 vssd1 vccd1 vccd1 _4992_/D sky130_fd_sc_hd__nor2_1
X_2525_ _2525_/A vssd1 vssd1 vccd1 vccd1 _5121_/D sky130_fd_sc_hd__clkbuf_1
X_5244_ _5446_/CLK _5244_/D vssd1 vssd1 vccd1 vccd1 _5580_/A sky130_fd_sc_hd__dfxtp_4
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _5351_/CLK _5175_/D vssd1 vssd1 vccd1 vccd1 _5175_/Q sky130_fd_sc_hd__dfxtp_2
X_4126_ _5342_/Q _5165_/Q _4126_/S vssd1 vssd1 vccd1 vccd1 _4127_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4057_ _5377_/Q hold70/A _4065_/S vssd1 vssd1 vccd1 vccd1 _4058_/A sky130_fd_sc_hd__mux2_1
X_3008_ _3134_/A _3008_/B vssd1 vssd1 vccd1 vccd1 _4832_/A sky130_fd_sc_hd__xnor2_4
XFILLER_52_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4959_ _5445_/Q _4959_/B _5446_/Q vssd1 vssd1 vccd1 vccd1 _4959_/X sky130_fd_sc_hd__or3b_1
XFILLER_137_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3290_ _3300_/A _3300_/B _3290_/C vssd1 vssd1 vccd1 vccd1 _3313_/B sky130_fd_sc_hd__nand3_1
XFILLER_3_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4813_ _4813_/A vssd1 vssd1 vccd1 vccd1 _5396_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4744_ _4744_/A _4744_/B vssd1 vssd1 vccd1 vccd1 _5355_/D sky130_fd_sc_hd__nor2_1
X_4675_ _3894_/B _4464_/C _4680_/B vssd1 vssd1 vccd1 vccd1 _4675_/Y sky130_fd_sc_hd__o21ai_1
X_3626_ _3643_/S vssd1 vssd1 vccd1 vccd1 _3626_/Y sky130_fd_sc_hd__inv_2
X_3557_ _4634_/A vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__clkbuf_4
X_3488_ _4042_/A _3472_/A _3486_/Y _3487_/Y vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__o211a_4
X_5227_ _5446_/CLK _5227_/D vssd1 vssd1 vccd1 vccd1 _5227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5158_ _5160_/CLK _5158_/D vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfxtp_1
X_4109_ _4109_/A _4109_/B vssd1 vssd1 vccd1 vccd1 _5159_/D sky130_fd_sc_hd__nor2_1
X_5089_ _5323_/CLK _5089_/D vssd1 vssd1 vccd1 vccd1 _5089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2790_ _2775_/X _2790_/B _3415_/A vssd1 vssd1 vccd1 vccd1 _4044_/A sky130_fd_sc_hd__nand3b_1
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4460_ _4353_/A _4457_/C _4459_/X _4416_/X vssd1 vssd1 vccd1 vccd1 _5253_/D sky130_fd_sc_hd__o211a_1
X_3411_ _3411_/A _3411_/B vssd1 vssd1 vccd1 vccd1 _3412_/A sky130_fd_sc_hd__nor2_1
X_4391_ _3654_/A _4383_/X _4390_/X _4378_/X vssd1 vssd1 vccd1 vccd1 _5234_/D sky130_fd_sc_hd__o211a_1
X_3342_ _3324_/A _3358_/A _3321_/A _3321_/B vssd1 vssd1 vccd1 vccd1 _3343_/B sky130_fd_sc_hd__a211o_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _3207_/B _3275_/B _3280_/A _3229_/B _3285_/B vssd1 vssd1 vccd1 vccd1 _3307_/B
+ sky130_fd_sc_hd__o311a_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5430_/CLK _5012_/D vssd1 vssd1 vccd1 vccd1 _5012_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2988_ _2985_/A _2987_/Y _2994_/A vssd1 vssd1 vccd1 vccd1 _2989_/B sky130_fd_sc_hd__mux2_1
X_4727_ _4727_/A _4727_/B vssd1 vssd1 vccd1 vccd1 _5334_/D sky130_fd_sc_hd__nor2_1
X_4658_ _5316_/Q _4657_/X _4662_/S vssd1 vssd1 vccd1 vccd1 _4659_/B sky130_fd_sc_hd__mux2_1
X_3609_ _5323_/Q vssd1 vssd1 vccd1 vccd1 _4504_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4589_ _4589_/A vssd1 vssd1 vccd1 vccd1 _4589_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3960_ _3960_/A vssd1 vssd1 vccd1 vccd1 _5092_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_16_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2911_ _2973_/A _2977_/A _2893_/X _2908_/X _2980_/A vssd1 vssd1 vccd1 vccd1 _2912_/B
+ sky130_fd_sc_hd__o221ai_4
X_3891_ _5000_/Q _3891_/B _3642_/A vssd1 vssd1 vccd1 vccd1 _3892_/A sky130_fd_sc_hd__nor3b_2
X_5630_ _5630_/A _2668_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__ebufn_8
X_2842_ _5021_/Q _5019_/Q _5020_/Q _5022_/Q _2860_/S _2833_/A vssd1 vssd1 vccd1 vccd1
+ _2842_/X sky130_fd_sc_hd__mux4_1
X_5561_ _5561_/A _2585_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[27] sky130_fd_sc_hd__ebufn_8
X_2773_ _5243_/Q _5231_/Q vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__nand2_1
X_4512_ _4512_/A vssd1 vssd1 vccd1 vccd1 _4515_/A sky130_fd_sc_hd__clkinv_2
Xhold104 hold126/X vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 _5063_/Q vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold115 hold96/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__clkbuf_1
Xhold137 _5369_/Q vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_4443_ _4434_/C _4438_/B _4355_/A vssd1 vssd1 vccd1 vccd1 _4443_/Y sky130_fd_sc_hd__o21ai_1
X_4374_ _5230_/Q _4362_/X _4373_/X _2750_/X vssd1 vssd1 vccd1 vccd1 _5230_/D sky130_fd_sc_hd__o211a_1
X_3325_ _3349_/A _3349_/B vssd1 vssd1 vccd1 vccd1 _3380_/A sky130_fd_sc_hd__and2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _3260_/A _3551_/C vssd1 vssd1 vccd1 vccd1 _3398_/A sky130_fd_sc_hd__nand2_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _3187_/A _5242_/Q vssd1 vssd1 vccd1 vccd1 _3187_/X sky130_fd_sc_hd__or2_1
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3110_ _3074_/A _5382_/Q _3076_/A _5313_/Q vssd1 vssd1 vccd1 vccd1 _3111_/B sky130_fd_sc_hd__a22o_1
X_4090_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4093_/A sky130_fd_sc_hd__buf_6
XFILLER_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3041_ _3041_/A vssd1 vssd1 vccd1 vccd1 _3084_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4992_ _5446_/CLK _4992_/D vssd1 vssd1 vccd1 vccd1 _4992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3943_ _3943_/A vssd1 vssd1 vccd1 vccd1 _3943_/X sky130_fd_sc_hd__clkbuf_2
X_3874_ _3874_/A vssd1 vssd1 vccd1 vccd1 _5070_/D sky130_fd_sc_hd__clkbuf_1
X_2825_ _2843_/S _2817_/X _2824_/X vssd1 vssd1 vccd1 vccd1 _2825_/Y sky130_fd_sc_hd__a21oi_1
X_5613_ _5613_/A _2647_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[9] sky130_fd_sc_hd__ebufn_8
X_2756_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4685_/A sky130_fd_sc_hd__clkbuf_4
X_5544_ _5544_/A _2693_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[10] sky130_fd_sc_hd__ebufn_8
X_2687_ _2689_/A vssd1 vssd1 vccd1 vccd1 _2687_/Y sky130_fd_sc_hd__inv_2
X_4426_ _5580_/A _4424_/X _4426_/S vssd1 vssd1 vccd1 vccd1 _4427_/B sky130_fd_sc_hd__mux2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _4357_/A _4450_/B vssd1 vssd1 vccd1 vccd1 _4357_/Y sky130_fd_sc_hd__nand2_1
X_3308_ _3354_/A _3354_/B vssd1 vssd1 vccd1 vccd1 _3308_/X sky130_fd_sc_hd__or2_1
X_4288_ _4287_/X _5213_/Q _4288_/S vssd1 vssd1 vccd1 vccd1 _4289_/A sky130_fd_sc_hd__mux2_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _3268_/A _3337_/A _3238_/X vssd1 vssd1 vccd1 vccd1 _3265_/B sky130_fd_sc_hd__a21bo_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_2
X_5476__66 vssd1 vssd1 vccd1 vccd1 _5476__66/HI _5553_/A sky130_fd_sc_hd__conb_1
XFILLER_18_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2610_ input1/X vssd1 vssd1 vccd1 vccd1 _2635_/A sky130_fd_sc_hd__buf_12
X_3590_ _5250_/Q vssd1 vssd1 vccd1 vccd1 _4449_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2541_ _5117_/Q _2541_/B vssd1 vssd1 vccd1 vccd1 _2546_/A sky130_fd_sc_hd__and2_1
X_5260_ _5435_/CLK _5260_/D vssd1 vssd1 vccd1 vccd1 _5260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4211_ _4210_/X _5192_/Q _4214_/S vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__mux2_1
X_5191_ _5369_/CLK _5191_/D vssd1 vssd1 vccd1 vccd1 _5191_/Q sky130_fd_sc_hd__dfxtp_1
X_4142_ hold138/X _5172_/Q _4148_/S vssd1 vssd1 vccd1 vccd1 _4143_/A sky130_fd_sc_hd__mux2_1
X_4073_ _3377_/A _4073_/B _4073_/C _4073_/D vssd1 vssd1 vccd1 vccd1 _4073_/X sky130_fd_sc_hd__and4b_1
XFILLER_49_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3024_ _3024_/A _3024_/B vssd1 vssd1 vccd1 vccd1 _4832_/B sky130_fd_sc_hd__xnor2_4
Xclkbuf_leaf_13_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5322_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5490__80 vssd1 vssd1 vccd1 vccd1 _5490__80/HI _5568_/A sky130_fd_sc_hd__conb_1
X_4975_ _4975_/A _4975_/B vssd1 vssd1 vccd1 vccd1 _4980_/B sky130_fd_sc_hd__nor2_1
XFILLER_24_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3926_ _5258_/Q _3919_/X _3897_/X _5080_/Q vssd1 vssd1 vccd1 vccd1 _3926_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3857_ _3857_/A vssd1 vssd1 vccd1 vccd1 _5062_/D sky130_fd_sc_hd__clkbuf_1
X_3788_ _3788_/A _3820_/A vssd1 vssd1 vccd1 vccd1 _3789_/A sky130_fd_sc_hd__and2_1
X_2808_ _5127_/Q _5128_/Q vssd1 vssd1 vccd1 vccd1 _3461_/A sky130_fd_sc_hd__or2_1
X_2739_ _2739_/A _2752_/B _2752_/C vssd1 vssd1 vccd1 vccd1 _2739_/Y sky130_fd_sc_hd__nor3_1
X_4409_ _4419_/A _4409_/B vssd1 vssd1 vccd1 vccd1 _4409_/X sky130_fd_sc_hd__or2_1
X_5389_ _5403_/Q _5389_/D vssd1 vssd1 vccd1 vccd1 _5389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4760_ _4765_/C _4760_/B vssd1 vssd1 vccd1 vccd1 _5360_/D sky130_fd_sc_hd__nor2_1
X_3711_ _4043_/A vssd1 vssd1 vccd1 vccd1 _3711_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4691_ _4692_/B _4588_/X _4690_/Y vssd1 vssd1 vccd1 vccd1 _5325_/D sky130_fd_sc_hd__o21a_1
X_3642_ _3642_/A _3642_/B vssd1 vssd1 vccd1 vccd1 _3642_/Y sky130_fd_sc_hd__nor2_1
X_5312_ _5313_/CLK _5312_/D vssd1 vssd1 vccd1 vccd1 _5312_/Q sky130_fd_sc_hd__dfxtp_1
X_3573_ _3572_/B _3571_/A _3569_/X vssd1 vssd1 vccd1 vccd1 _3574_/B sky130_fd_sc_hd__o21ai_1
XFILLER_5_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2524_ _5587_/A _2527_/B _2548_/C vssd1 vssd1 vccd1 vccd1 _2525_/A sky130_fd_sc_hd__and3_1
X_5243_ _5445_/CLK _5243_/D vssd1 vssd1 vccd1 vccd1 _5243_/Q sky130_fd_sc_hd__dfxtp_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ _5351_/CLK _5174_/D vssd1 vssd1 vccd1 vccd1 _5174_/Q sky130_fd_sc_hd__dfxtp_2
X_4125_ _4125_/A vssd1 vssd1 vccd1 vccd1 _5164_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4056_ _4071_/S vssd1 vssd1 vccd1 vccd1 _4065_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_43_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3007_ _3041_/A _3013_/B _3004_/Y _3006_/Y vssd1 vssd1 vccd1 vccd1 _3008_/B sky130_fd_sc_hd__o22a_1
XFILLER_24_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4958_ _5445_/Q _4959_/B vssd1 vssd1 vccd1 vccd1 _4958_/Y sky130_fd_sc_hd__nand2_1
X_4889_ _5414_/Q _4888_/C _5415_/Q vssd1 vssd1 vccd1 vccd1 _4889_/Y sky130_fd_sc_hd__a21oi_1
X_3909_ _3956_/S vssd1 vssd1 vccd1 vccd1 _3909_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5460__50 vssd1 vssd1 vccd1 vccd1 _5460__50/HI _5537_/A sky130_fd_sc_hd__conb_1
X_4812_ _4834_/A _5396_/Q _4812_/S vssd1 vssd1 vccd1 vccd1 _4813_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4743_ _5355_/Q _4742_/X _5371_/D vssd1 vssd1 vccd1 vccd1 _4744_/B sky130_fd_sc_hd__a21oi_1
X_4674_ _4674_/A _4464_/C vssd1 vssd1 vccd1 vccd1 _4680_/B sky130_fd_sc_hd__or2b_1
X_5527__117 vssd1 vssd1 vccd1 vccd1 _5527__117/HI _5527__117/LO sky130_fd_sc_hd__conb_1
X_3625_ _4708_/A _3946_/A _3625_/C vssd1 vssd1 vccd1 vccd1 _3643_/S sky130_fd_sc_hd__or3_2
X_3556_ _3556_/A vssd1 vssd1 vccd1 vccd1 _4987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5226_ _5328_/CLK _5226_/D vssd1 vssd1 vccd1 vccd1 _5579_/A sky130_fd_sc_hd__dfxtp_1
X_3487_ _4042_/A _3472_/A _3489_/A vssd1 vssd1 vccd1 vccd1 _3487_/Y sky130_fd_sc_hd__a21oi_1
X_5157_ _5313_/CLK _5157_/D vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfxtp_1
X_4108_ hold43/A _4106_/A _2766_/A vssd1 vssd1 vccd1 vccd1 _4109_/B sky130_fd_sc_hd__o21ai_1
X_5088_ _5435_/CLK _5088_/D vssd1 vssd1 vccd1 vccd1 _5088_/Q sky130_fd_sc_hd__dfxtp_1
X_4039_ _4038_/A _2823_/Y _4022_/B _4038_/Y vssd1 vssd1 vccd1 vccd1 _4039_/X sky130_fd_sc_hd__o211a_1
XFILLER_24_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3410_ _3388_/A _3388_/B _3314_/X vssd1 vssd1 vccd1 vccd1 _3413_/A sky130_fd_sc_hd__a21o_1
X_4390_ _4400_/A _4390_/B vssd1 vssd1 vccd1 vccd1 _4390_/X sky130_fd_sc_hd__or2_1
X_3341_ _3344_/A _3341_/B vssd1 vssd1 vccd1 vccd1 _3372_/A sky130_fd_sc_hd__nor2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _5442_/Q _3272_/B vssd1 vssd1 vccd1 vccd1 _3280_/A sky130_fd_sc_hd__nor2_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5011_ _5430_/CLK _5011_/D vssd1 vssd1 vccd1 vccd1 _5011_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2987_ _2987_/A _2987_/B vssd1 vssd1 vccd1 vccd1 _2987_/Y sky130_fd_sc_hd__xnor2_1
X_4003__10 _4002__9/A vssd1 vssd1 vccd1 vccd1 _5117_/CLK sky130_fd_sc_hd__inv_2
X_4726_ _5334_/Q _4724_/A _4710_/B vssd1 vssd1 vccd1 vccd1 _4727_/B sky130_fd_sc_hd__o21ai_1
X_4657_ _5298_/Q _5268_/Q _4661_/S vssd1 vssd1 vccd1 vccd1 _4657_/X sky130_fd_sc_hd__mux2_1
X_3608_ _4999_/Q _3602_/X _3606_/X _3608_/B2 vssd1 vssd1 vccd1 vccd1 _4999_/D sky130_fd_sc_hd__a22o_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4588_ _4591_/A vssd1 vssd1 vccd1 vccd1 _4588_/X sky130_fd_sc_hd__clkbuf_2
X_3539_ _3682_/B _3682_/C _3539_/C vssd1 vssd1 vccd1 vccd1 _3539_/X sky130_fd_sc_hd__and3_1
X_5209_ _5339_/CLK _5209_/D vssd1 vssd1 vccd1 vccd1 _5209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2910_ _2910_/A vssd1 vssd1 vccd1 vccd1 _2980_/A sky130_fd_sc_hd__clkbuf_2
X_3890_ _5324_/Q vssd1 vssd1 vccd1 vccd1 _4692_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2841_ _2839_/X _5016_/Q _5015_/Q _5018_/Q _2833_/A _2860_/S vssd1 vssd1 vccd1 vccd1
+ _2841_/X sky130_fd_sc_hd__mux4_1
X_5560_ _5560_/A _2584_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[26] sky130_fd_sc_hd__ebufn_8
X_2772_ _4829_/S _5419_/Q vssd1 vssd1 vccd1 vccd1 _4959_/B sky130_fd_sc_hd__nand2_2
X_4511_ _5271_/Q _5272_/Q _4514_/B vssd1 vssd1 vccd1 vccd1 _4512_/A sky130_fd_sc_hd__or3_1
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold127/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold116 hold99/X vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__clkbuf_2
X_4442_ _5247_/Q _4438_/B _4441_/X _4093_/A vssd1 vssd1 vccd1 vccd1 _5247_/D sky130_fd_sc_hd__a211o_1
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold138 _5349_/Q vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_4373_ _4381_/A _4373_/B vssd1 vssd1 vccd1 vccd1 _4373_/X sky130_fd_sc_hd__or2_1
X_3324_ _3324_/A _3334_/A vssd1 vssd1 vccd1 vccd1 _3349_/B sky130_fd_sc_hd__or2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _4993_/Q vssd1 vssd1 vccd1 vccd1 _3551_/C sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _4835_/B vssd1 vssd1 vccd1 vccd1 _3186_/X sky130_fd_sc_hd__buf_2
XFILLER_39_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_wb_clk_i clkbuf_2_3_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_50_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4709_ _4720_/C vssd1 vssd1 vccd1 vccd1 _4710_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3040_ _3040_/A _3040_/B vssd1 vssd1 vccd1 vccd1 _3040_/Y sky130_fd_sc_hd__xnor2_1
X_4991_ _5439_/CLK _4991_/D vssd1 vssd1 vccd1 vccd1 _4991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _3946_/A _3942_/B vssd1 vssd1 vccd1 vccd1 _3943_/A sky130_fd_sc_hd__or2_1
X_3873_ hold13/A _4833_/B _3873_/S vssd1 vssd1 vccd1 vccd1 _3874_/A sky130_fd_sc_hd__mux2_1
X_5612_ _5612_/A _2646_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[8] sky130_fd_sc_hd__ebufn_8
X_2824_ _2823_/Y _2838_/A _2824_/S vssd1 vssd1 vccd1 vccd1 _2824_/X sky130_fd_sc_hd__mux2_1
X_5543_ _5543_/A _2694_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[9] sky130_fd_sc_hd__ebufn_8
XFILLER_8_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2755_ _2760_/A _2768_/A vssd1 vssd1 vccd1 vccd1 _2755_/X sky130_fd_sc_hd__or2b_1
X_2686_ _2689_/A vssd1 vssd1 vccd1 vccd1 _2686_/Y sky130_fd_sc_hd__inv_2
X_4425_ _4355_/A _3674_/B _4363_/C _4739_/A vssd1 vssd1 vccd1 vccd1 _4426_/S sky130_fd_sc_hd__o211a_1
X_4356_ _4432_/A _4434_/B _4450_/B vssd1 vssd1 vccd1 vccd1 _4356_/X sky130_fd_sc_hd__o21a_1
X_3307_ _3309_/A _3307_/B vssd1 vssd1 vccd1 vccd1 _3354_/B sky130_fd_sc_hd__xnor2_1
XFILLER_48_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ _5209_/Q _4275_/X _4286_/X vssd1 vssd1 vccd1 vccd1 _4287_/X sky130_fd_sc_hd__a21o_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _3238_/A _3233_/B vssd1 vssd1 vccd1 vccd1 _3238_/X sky130_fd_sc_hd__or2b_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3169_ _3654_/A _3169_/B vssd1 vssd1 vccd1 vccd1 _4835_/A sky130_fd_sc_hd__xor2_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2540_ _5116_/Q _2734_/A _2554_/A vssd1 vssd1 vccd1 vccd1 _2541_/B sky130_fd_sc_hd__and3_1
X_4210_ _5416_/Q _5367_/Q _4216_/S vssd1 vssd1 vccd1 vccd1 _4210_/X sky130_fd_sc_hd__mux2_1
X_5190_ _5369_/CLK _5190_/D vssd1 vssd1 vccd1 vccd1 _5190_/Q sky130_fd_sc_hd__dfxtp_1
X_4141_ _4141_/A vssd1 vssd1 vccd1 vccd1 _5171_/D sky130_fd_sc_hd__clkbuf_1
X_4072_ _4072_/A vssd1 vssd1 vccd1 vccd1 _5147_/D sky130_fd_sc_hd__clkbuf_1
X_3023_ _3023_/A _3023_/B vssd1 vssd1 vccd1 vccd1 _3024_/B sky130_fd_sc_hd__xnor2_2
XFILLER_36_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4974_ _4975_/A _4975_/B vssd1 vssd1 vccd1 vccd1 _4982_/B sky130_fd_sc_hd__or2_1
X_3925_ _5083_/Q _3909_/X _3924_/X vssd1 vssd1 vccd1 vccd1 _5083_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3856_ _5062_/Q _2918_/X _5133_/D vssd1 vssd1 vccd1 vccd1 _3857_/A sky130_fd_sc_hd__mux2_1
XFILLER_20_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2807_ _5129_/Q vssd1 vssd1 vccd1 vccd1 _3464_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3787_ _3805_/C vssd1 vssd1 vccd1 vccd1 _3820_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2738_ _5118_/Q _5111_/Q _5110_/Q _5113_/Q vssd1 vssd1 vccd1 vccd1 _2752_/C sky130_fd_sc_hd__or4b_1
X_2669_ _2671_/A vssd1 vssd1 vccd1 vccd1 _2669_/Y sky130_fd_sc_hd__inv_2
X_4408_ _5202_/Q _5172_/Q _4418_/S vssd1 vssd1 vccd1 vccd1 _4409_/B sky130_fd_sc_hd__mux2_1
X_5388_ _5403_/Q _5388_/D vssd1 vssd1 vccd1 vccd1 _5388_/Q sky130_fd_sc_hd__dfxtp_1
X_4339_ _5577_/A _4338_/X _4347_/S vssd1 vssd1 vccd1 vccd1 _4340_/B sky130_fd_sc_hd__mux2_1
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3710_ _3720_/B _4043_/A _3736_/A vssd1 vssd1 vccd1 vccd1 _3710_/X sky130_fd_sc_hd__and3_1
X_4690_ _4588_/X _4689_/X _4094_/X vssd1 vssd1 vccd1 vccd1 _4690_/Y sky130_fd_sc_hd__a21oi_1
X_3641_ _4587_/A _3641_/B vssd1 vssd1 vccd1 vccd1 _3642_/B sky130_fd_sc_hd__and2b_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3572_ _3572_/A _3572_/B _3575_/B vssd1 vssd1 vccd1 vccd1 _3574_/A sky130_fd_sc_hd__and3_1
X_5311_ _5328_/CLK _5311_/D vssd1 vssd1 vccd1 vccd1 _5311_/Q sky130_fd_sc_hd__dfxtp_1
X_2523_ _2768_/A _5586_/A vssd1 vssd1 vccd1 vccd1 _2548_/C sky130_fd_sc_hd__nor2_2
XFILLER_5_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5242_ _5445_/CLK _5242_/D vssd1 vssd1 vccd1 vccd1 _5242_/Q sky130_fd_sc_hd__dfxtp_1
X_5173_ _5351_/CLK _5173_/D vssd1 vssd1 vccd1 vccd1 _5173_/Q sky130_fd_sc_hd__dfxtp_2
X_4124_ _5341_/Q _5164_/Q _4126_/S vssd1 vssd1 vccd1 vccd1 _4125_/A sky130_fd_sc_hd__mux2_1
Xinput1 active vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_6
X_4055_ _4055_/A vssd1 vssd1 vccd1 vccd1 _5139_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3006_ _3041_/A _3013_/C vssd1 vssd1 vccd1 vccd1 _3006_/Y sky130_fd_sc_hd__nand2_1
X_4957_ _4842_/X _4959_/B input20/X vssd1 vssd1 vccd1 vccd1 _5444_/D sky130_fd_sc_hd__a21boi_1
X_4888_ _5414_/Q _5415_/Q _4888_/C vssd1 vssd1 vccd1 vccd1 _4893_/B sky130_fd_sc_hd__and3_1
X_3908_ _3908_/A vssd1 vssd1 vccd1 vccd1 _5080_/D sky130_fd_sc_hd__clkbuf_1
X_3839_ _3841_/B _3847_/C _3854_/A vssd1 vssd1 vccd1 vccd1 _3839_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_20_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4811_ _4811_/A vssd1 vssd1 vccd1 vccd1 _5395_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4742_ _4762_/A vssd1 vssd1 vccd1 vccd1 _4742_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4673_ _4673_/A vssd1 vssd1 vccd1 vccd1 _5319_/D sky130_fd_sc_hd__clkbuf_1
X_3624_ _3912_/A _3623_/X _5254_/Q vssd1 vssd1 vccd1 vccd1 _3625_/C sky130_fd_sc_hd__o21ai_1
X_3555_ _3377_/A _3569_/A vssd1 vssd1 vccd1 vccd1 _3556_/A sky130_fd_sc_hd__and2b_1
X_3486_ _3467_/X _3473_/Y _3485_/X vssd1 vssd1 vccd1 vccd1 _3486_/Y sky130_fd_sc_hd__o21ai_1
X_5225_ _5328_/CLK _5225_/D vssd1 vssd1 vccd1 vccd1 _5578_/A sky130_fd_sc_hd__dfxtp_1
X_5156_ _5313_/CLK _5156_/D vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4107_ hold43/A hold46/A _4107_/C vssd1 vssd1 vccd1 vccd1 _4109_/A sky130_fd_sc_hd__and3_1
X_5087_ _5435_/CLK _5087_/D vssd1 vssd1 vccd1 vccd1 _5087_/Q sky130_fd_sc_hd__dfxtp_1
X_4038_ _4038_/A _4038_/B vssd1 vssd1 vccd1 vccd1 _4038_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5510__100 vssd1 vssd1 vccd1 vccd1 _5510__100/HI _5613_/A sky130_fd_sc_hd__conb_1
XFILLER_4_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5506__96 vssd1 vssd1 vccd1 vccd1 _5506__96/HI _5609_/A sky130_fd_sc_hd__conb_1
XFILLER_0_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3340_ _3352_/S _3340_/B vssd1 vssd1 vccd1 vccd1 _3340_/Y sky130_fd_sc_hd__nand2_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3251_/A _3250_/A _3249_/X vssd1 vssd1 vccd1 vccd1 _3272_/B sky130_fd_sc_hd__o21a_1
X_5010_ _5444_/CLK _5010_/D vssd1 vssd1 vccd1 vccd1 _5010_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2986_ _2961_/A _2961_/B _2962_/Y vssd1 vssd1 vccd1 vccd1 _2987_/B sky130_fd_sc_hd__a21o_1
XFILLER_30_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4725_ _5333_/Q _5334_/Q _4725_/C vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__and3_1
X_4656_ _4656_/A vssd1 vssd1 vccd1 vccd1 _5315_/D sky130_fd_sc_hd__clkbuf_1
X_3607_ _4998_/Q _3602_/X _3606_/X _3607_/B2 vssd1 vssd1 vccd1 vccd1 _4998_/D sky130_fd_sc_hd__a22o_1
X_4587_ _4587_/A _4587_/B _4587_/C vssd1 vssd1 vccd1 vccd1 _4591_/A sky130_fd_sc_hd__and3_1
X_3538_ _3530_/X _3535_/X _3537_/X _5174_/Q vssd1 vssd1 vccd1 vccd1 _3539_/C sky130_fd_sc_hd__a22o_1
X_3469_ _2810_/X _2813_/Y _3468_/X vssd1 vssd1 vccd1 vccd1 _3469_/X sky130_fd_sc_hd__a21o_1
X_5208_ _5369_/CLK _5208_/D vssd1 vssd1 vccd1 vccd1 _5208_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0_0__1653_ clkbuf_0__1653_/X vssd1 vssd1 vccd1 vccd1 _4002__9/A sky130_fd_sc_hd__clkbuf_2
X_5139_ _5313_/CLK _5139_/D vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5335_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2840_ _2840_/A vssd1 vssd1 vccd1 vccd1 _2860_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_31_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2771_ _5403_/Q vssd1 vssd1 vccd1 vccd1 _4829_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_8_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4510_ _5271_/Q _4514_/B _4509_/X vssd1 vssd1 vccd1 vccd1 _5271_/D sky130_fd_sc_hd__a21bo_1
Xhold106 hold130/X vssd1 vssd1 vccd1 vccd1 hold107/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 hold98/X vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__clkbuf_1
X_4441_ _4434_/C _3674_/B _4438_/B vssd1 vssd1 vccd1 vccd1 _4441_/X sky130_fd_sc_hd__o21ba_1
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold139 _5335_/Q vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__clkdlybuf4s25_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ input8/X _5163_/Q _4380_/S vssd1 vssd1 vccd1 vccd1 _4373_/B sky130_fd_sc_hd__mux2_1
X_3323_ _3328_/A _3559_/B vssd1 vssd1 vccd1 vccd1 _3334_/A sky130_fd_sc_hd__nand2_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5497__87 vssd1 vssd1 vccd1 vccd1 _5497__87/HI _5596_/A sky130_fd_sc_hd__conb_1
XFILLER_58_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3254_ _3260_/A _4993_/Q vssd1 vssd1 vccd1 vccd1 _3438_/B sky130_fd_sc_hd__or2_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _3654_/A _3185_/B vssd1 vssd1 vccd1 vccd1 _4835_/B sky130_fd_sc_hd__xnor2_1
XFILLER_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2969_ _3029_/A vssd1 vssd1 vccd1 vccd1 _3108_/A sky130_fd_sc_hd__clkbuf_1
X_4708_ _4708_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _4720_/C sky130_fd_sc_hd__nor2_1
X_4639_ _5294_/Q _5264_/Q _4639_/S vssd1 vssd1 vccd1 vccd1 _4639_/X sky130_fd_sc_hd__mux2_1
XFILLER_49_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4990_ _5335_/CLK _4990_/D vssd1 vssd1 vccd1 vccd1 _4990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3941_ hold133/X _3932_/X _3904_/C _3940_/X vssd1 vssd1 vccd1 vccd1 _5088_/D sky130_fd_sc_hd__a31o_1
X_3872_ _3872_/A vssd1 vssd1 vccd1 vccd1 _5069_/D sky130_fd_sc_hd__clkbuf_1
X_5611_ _5611_/A _2645_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[7] sky130_fd_sc_hd__ebufn_8
X_2823_ _3462_/B _2823_/B vssd1 vssd1 vccd1 vccd1 _2823_/Y sky130_fd_sc_hd__nand2_1
X_5542_ _5542_/A _2695_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[8] sky130_fd_sc_hd__ebufn_8
X_2754_ _5150_/Q vssd1 vssd1 vccd1 vccd1 _2760_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2685_ _2689_/A vssd1 vssd1 vccd1 vccd1 _2685_/Y sky130_fd_sc_hd__inv_2
X_4424_ _4432_/A _3528_/A _4353_/X _3511_/Y _4363_/B vssd1 vssd1 vccd1 vccd1 _4424_/X
+ sky130_fd_sc_hd__a311o_1
X_4355_ _4355_/A _5247_/Q _4355_/C vssd1 vssd1 vccd1 vccd1 _4450_/B sky130_fd_sc_hd__and3_1
X_3306_ _3306_/A _3306_/B vssd1 vssd1 vccd1 vccd1 _3354_/A sky130_fd_sc_hd__nor2_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _5163_/Q _4285_/X _4276_/X _5189_/Q vssd1 vssd1 vccd1 vccd1 _4286_/X sky130_fd_sc_hd__a22o_1
X_3237_ _3336_/A _3349_/A vssd1 vssd1 vccd1 vccd1 _3337_/A sky130_fd_sc_hd__nor2_2
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3168_ _3649_/A _3181_/B _3166_/Y _3167_/Y vssd1 vssd1 vccd1 vccd1 _3169_/B sky130_fd_sc_hd__a31o_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3099_ _3099_/A vssd1 vssd1 vccd1 vccd1 _3100_/B sky130_fd_sc_hd__inv_2
XFILLER_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4140_ _5348_/Q _5171_/Q _4148_/S vssd1 vssd1 vccd1 vccd1 _4141_/A sky130_fd_sc_hd__mux2_1
X_4071_ _5384_/Q hold82/A _4071_/S vssd1 vssd1 vccd1 vccd1 _4072_/A sky130_fd_sc_hd__mux2_1
X_5467__57 vssd1 vssd1 vccd1 vccd1 _5467__57/HI _5544_/A sky130_fd_sc_hd__conb_1
X_3022_ _3090_/A _3021_/A _3067_/B vssd1 vssd1 vccd1 vccd1 _3023_/B sky130_fd_sc_hd__a21boi_1
XFILLER_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _2990_/X _4965_/Y _4972_/X _4902_/X vssd1 vssd1 vccd1 vccd1 _5450_/D sky130_fd_sc_hd__o211a_1
X_3924_ _5283_/Q _3910_/X _3911_/X _3923_/X vssd1 vssd1 vccd1 vccd1 _3924_/X sky130_fd_sc_hd__a211o_1
XFILLER_32_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3855_ _3855_/A vssd1 vssd1 vccd1 vccd1 _5061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2806_ _5027_/Q _5028_/Q _2869_/A vssd1 vssd1 vccd1 vccd1 _2806_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0__1653_ _4000_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__1653_/X sky130_fd_sc_hd__clkbuf_16
X_3786_ _2713_/B _2728_/X _2764_/X _3785_/Y _3698_/A vssd1 vssd1 vccd1 vccd1 _3805_/C
+ sky130_fd_sc_hd__o41a_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5305_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_2737_ _2729_/C _5116_/Q _2737_/C _2737_/D vssd1 vssd1 vccd1 vccd1 _2759_/A sky130_fd_sc_hd__and4bb_1
X_2668_ _2671_/A vssd1 vssd1 vccd1 vccd1 _2668_/Y sky130_fd_sc_hd__inv_2
X_4407_ _3648_/A _4402_/X _4406_/X _4397_/X vssd1 vssd1 vccd1 vccd1 _5238_/D sky130_fd_sc_hd__o211a_1
X_2599_ _2603_/A vssd1 vssd1 vccd1 vccd1 _2599_/Y sky130_fd_sc_hd__inv_2
X_5387_ _5403_/Q _5387_/D vssd1 vssd1 vccd1 vccd1 _5387_/Q sky130_fd_sc_hd__dfxtp_1
X_4338_ _5268_/Q _3919_/A _3943_/X _5090_/Q _3947_/X vssd1 vssd1 vccd1 vccd1 _4338_/X
+ sky130_fd_sc_hd__a221o_1
X_4269_ _4292_/A vssd1 vssd1 vccd1 vccd1 _4288_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5481__71 vssd1 vssd1 vccd1 vccd1 _5481__71/HI _5558_/A sky130_fd_sc_hd__conb_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3640_ _4594_/A vssd1 vssd1 vccd1 vccd1 _4587_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3571_ _3571_/A _3571_/B vssd1 vssd1 vccd1 vccd1 _4991_/D sky130_fd_sc_hd__nor2_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5310_ _5436_/CLK _5310_/D vssd1 vssd1 vccd1 vccd1 _5310_/Q sky130_fd_sc_hd__dfxtp_1
X_2522_ _5038_/Q vssd1 vssd1 vccd1 vccd1 _2768_/A sky130_fd_sc_hd__clkbuf_2
X_5241_ _5445_/CLK _5241_/D vssd1 vssd1 vccd1 vccd1 _5241_/Q sky130_fd_sc_hd__dfxtp_1
X_5172_ _5351_/CLK _5172_/D vssd1 vssd1 vccd1 vccd1 _5172_/Q sky130_fd_sc_hd__dfxtp_2
X_4123_ _4123_/A vssd1 vssd1 vccd1 vccd1 _5163_/D sky130_fd_sc_hd__clkbuf_1
Xinput2 io_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_6
X_4054_ _5376_/Q hold79/A _4054_/S vssd1 vssd1 vccd1 vccd1 _4055_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3005_ _3005_/A _3065_/A vssd1 vssd1 vccd1 vccd1 _3013_/C sky130_fd_sc_hd__nand2_1
XFILLER_36_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ _5443_/Q _4954_/C _4955_/Y vssd1 vssd1 vccd1 vccd1 _5443_/D sky130_fd_sc_hd__o21a_1
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3907_ _5080_/Q _3906_/X _3956_/S vssd1 vssd1 vccd1 vccd1 _3908_/A sky130_fd_sc_hd__mux2_1
X_4887_ _5382_/D _4884_/X _4886_/Y _4882_/X vssd1 vssd1 vccd1 vccd1 _5414_/D sky130_fd_sc_hd__o211a_1
XFILLER_137_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3838_ _3838_/A vssd1 vssd1 vccd1 vccd1 _3854_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3769_ _3769_/A0 _3769_/A1 _3773_/S vssd1 vssd1 vccd1 vccd1 _3769_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5439_ _5439_/CLK _5439_/D vssd1 vssd1 vccd1 vccd1 _5439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4810_ _4833_/B _5395_/Q _4812_/S vssd1 vssd1 vccd1 vccd1 _4811_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _5109_/Q _4203_/A vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__or2b_1
XFILLER_21_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4672_ _4685_/A _4672_/B vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__or2_1
X_3623_ _5301_/Q _3912_/B _3895_/A vssd1 vssd1 vccd1 vccd1 _3623_/X sky130_fd_sc_hd__o21a_1
X_3554_ _4708_/A _3829_/C vssd1 vssd1 vccd1 vccd1 _3569_/A sky130_fd_sc_hd__nor2_2
XFILLER_6_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3485_ _4038_/B _3479_/Y _3484_/Y _3470_/Y vssd1 vssd1 vccd1 vccd1 _3485_/X sky130_fd_sc_hd__a211o_1
X_5224_ _5328_/CLK _5224_/D vssd1 vssd1 vccd1 vccd1 _5577_/A sky130_fd_sc_hd__dfxtp_1
X_5155_ _5160_/CLK _5155_/D vssd1 vssd1 vccd1 vccd1 _5155_/Q sky130_fd_sc_hd__dfxtp_4
X_4106_ _4106_/A _4106_/B vssd1 vssd1 vccd1 vccd1 _5158_/D sky130_fd_sc_hd__nor2_1
X_5086_ _5323_/CLK _5086_/D vssd1 vssd1 vccd1 vccd1 _5086_/Q sky130_fd_sc_hd__dfxtp_1
X_4037_ _2854_/Y _4030_/Y _4035_/X _4036_/Y _4043_/A vssd1 vssd1 vccd1 vccd1 _5130_/D
+ sky130_fd_sc_hd__a221oi_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4939_ _4939_/A vssd1 vssd1 vccd1 vccd1 _5434_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3270_ _3251_/A _3250_/A _3249_/X _5442_/Q vssd1 vssd1 vccd1 vccd1 _3275_/B sky130_fd_sc_hd__o211a_1
XFILLER_3_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5533__123 vssd1 vssd1 vccd1 vccd1 _5533__123/HI _5533__123/LO sky130_fd_sc_hd__conb_1
XFILLER_21_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4724_ _4724_/A _4724_/B vssd1 vssd1 vccd1 vccd1 _5333_/D sky130_fd_sc_hd__nor2_1
X_2985_ _2985_/A _2984_/Y vssd1 vssd1 vccd1 vccd1 _2987_/A sky130_fd_sc_hd__or2b_1
XFILLER_30_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4655_ _4655_/A _4655_/B vssd1 vssd1 vccd1 vccd1 _4656_/A sky130_fd_sc_hd__and2_1
X_3606_ _3606_/A _3726_/A _3729_/B vssd1 vssd1 vccd1 vccd1 _3606_/X sky130_fd_sc_hd__and3_1
X_4586_ _4586_/A _5327_/Q _4586_/C _4586_/D vssd1 vssd1 vccd1 vccd1 _4586_/X sky130_fd_sc_hd__and4_1
X_3537_ _4285_/A vssd1 vssd1 vccd1 vccd1 _3537_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3468_ _4034_/A _2824_/S _2806_/X vssd1 vssd1 vccd1 vccd1 _3468_/X sky130_fd_sc_hd__o21a_1
X_3399_ _3348_/X _3349_/A _3398_/X vssd1 vssd1 vccd1 vccd1 _3399_/Y sky130_fd_sc_hd__a21oi_1
X_5207_ _5245_/CLK _5207_/D vssd1 vssd1 vccd1 vccd1 _5207_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0__1652_ clkbuf_0__1652_/X vssd1 vssd1 vccd1 vccd1 _3999__7/A sky130_fd_sc_hd__clkbuf_2
X_5138_ _5313_/CLK _5138_/D vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5069_ _5077_/CLK _5069_/D vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5517__107 vssd1 vssd1 vccd1 vccd1 _5517__107/HI _5633_/A sky130_fd_sc_hd__conb_1
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2770_ _5385_/Q vssd1 vssd1 vccd1 vccd1 _2889_/B sky130_fd_sc_hd__clkbuf_4
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold131/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_8_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4440_ _4450_/A _4438_/Y _4439_/Y vssd1 vssd1 vccd1 vccd1 _5246_/D sky130_fd_sc_hd__a21oi_1
Xhold118 _5153_/Q vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_4371_ _5229_/Q _4362_/X _4370_/X _2750_/X vssd1 vssd1 vccd1 vccd1 _5229_/D sky130_fd_sc_hd__o211a_1
X_3322_ _4989_/Q vssd1 vssd1 vccd1 vccd1 _3324_/A sky130_fd_sc_hd__inv_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3260_/A vssd1 vssd1 vccd1 vccd1 _3572_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3184_ _3646_/A _3181_/X _3646_/C _3183_/Y vssd1 vssd1 vccd1 vccd1 _3185_/B sky130_fd_sc_hd__o31a_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2968_ _5238_/Q vssd1 vssd1 vccd1 vccd1 _3051_/A sky130_fd_sc_hd__clkbuf_2
X_4707_ _4707_/A _4707_/B _4707_/C vssd1 vssd1 vccd1 vccd1 _4827_/B sky130_fd_sc_hd__nor3_1
X_4638_ _4638_/A vssd1 vssd1 vccd1 vccd1 _5311_/D sky130_fd_sc_hd__clkbuf_1
X_2899_ _2953_/B _2953_/C vssd1 vssd1 vccd1 vccd1 _4975_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4569_ _5290_/Q _4566_/X _4568_/X _4558_/X vssd1 vssd1 vccd1 vccd1 _5294_/D sky130_fd_sc_hd__o211a_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3940_ _5088_/Q _3939_/X _3959_/S vssd1 vssd1 vccd1 vccd1 _3940_/X sky130_fd_sc_hd__mux2_1
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3871_ hold22/A _4832_/C _3873_/S vssd1 vssd1 vccd1 vccd1 _3872_/A sky130_fd_sc_hd__mux2_1
X_2822_ _2838_/A _2822_/B vssd1 vssd1 vccd1 vccd1 _2823_/B sky130_fd_sc_hd__nand2_1
X_5610_ _5610_/A _2644_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[6] sky130_fd_sc_hd__ebufn_8
X_5541_ _5541_/A _2696_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[7] sky130_fd_sc_hd__ebufn_8
X_2753_ _2753_/A _2753_/B vssd1 vssd1 vccd1 vccd1 _2753_/Y sky130_fd_sc_hd__nand2_1
X_2684_ _2690_/A vssd1 vssd1 vccd1 vccd1 _2689_/A sky130_fd_sc_hd__buf_2
X_4423_ _2991_/A _4402_/A _4422_/X _4416_/X vssd1 vssd1 vccd1 vccd1 _5243_/D sky130_fd_sc_hd__o211a_1
X_4354_ _4449_/C vssd1 vssd1 vccd1 vccd1 _4357_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3305_ _3396_/A _3305_/B vssd1 vssd1 vccd1 vccd1 _3306_/B sky130_fd_sc_hd__and2_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _4285_/A vssd1 vssd1 vccd1 vccd1 _4285_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3236_ _4989_/Q _3559_/B _3328_/A vssd1 vssd1 vccd1 vccd1 _3349_/A sky130_fd_sc_hd__o21a_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3167_ _3649_/A _3181_/A vssd1 vssd1 vccd1 vccd1 _3167_/Y sky130_fd_sc_hd__nor2_1
X_3098_ _3097_/A _3097_/B _3097_/C vssd1 vssd1 vccd1 vccd1 _3099_/A sky130_fd_sc_hd__o21a_1
XFILLER_27_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4070_ _4070_/A vssd1 vssd1 vccd1 vccd1 _5146_/D sky130_fd_sc_hd__clkbuf_1
X_3021_ _3021_/A _3021_/B vssd1 vssd1 vccd1 vccd1 _3067_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4972_ _4965_/A _4965_/B _5603_/A vssd1 vssd1 vccd1 vccd1 _4972_/X sky130_fd_sc_hd__a21o_1
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3923_ _5257_/Q _3915_/X _3897_/X _5079_/Q vssd1 vssd1 vccd1 vccd1 _3923_/X sky130_fd_sc_hd__a22o_1
X_3854_ _3854_/A _3854_/B vssd1 vssd1 vccd1 vccd1 _3855_/A sky130_fd_sc_hd__and2_1
XFILLER_137_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2805_ _2824_/S _2813_/B vssd1 vssd1 vccd1 vccd1 _2826_/A sky130_fd_sc_hd__or2_1
Xclkbuf_0__1652_ _3994_/X vssd1 vssd1 vccd1 vccd1 clkbuf_0__1652_/X sky130_fd_sc_hd__clkbuf_16
X_3785_ _5038_/Q _4075_/A _2753_/Y _2759_/X vssd1 vssd1 vccd1 vccd1 _3785_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2736_ _5117_/Q _2736_/B _2739_/A _5110_/Q vssd1 vssd1 vccd1 vccd1 _2737_/D sky130_fd_sc_hd__and4_1
X_2667_ _2671_/A vssd1 vssd1 vccd1 vccd1 _2667_/Y sky130_fd_sc_hd__inv_2
X_4406_ _4419_/A _4406_/B vssd1 vssd1 vccd1 vccd1 _4406_/X sky130_fd_sc_hd__or2_1
X_2598_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2603_/A sky130_fd_sc_hd__clkbuf_2
X_5386_ _5403_/Q _5386_/D vssd1 vssd1 vccd1 vccd1 _5386_/Q sky130_fd_sc_hd__dfxtp_1
X_4337_ _4327_/X _4335_/Y _4336_/Y vssd1 vssd1 vccd1 vccd1 _5223_/D sky130_fd_sc_hd__o21ai_1
X_4268_ _5185_/Q _3682_/D _4264_/X _5009_/Q vssd1 vssd1 vccd1 vccd1 _4268_/X sky130_fd_sc_hd__a22o_1
X_3219_ _3829_/B _3277_/B _5439_/Q vssd1 vssd1 vccd1 vccd1 _3221_/B sky130_fd_sc_hd__o21a_1
XFILLER_27_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4199_ _5413_/Q _5364_/Q _4199_/S vssd1 vssd1 vccd1 vccd1 _4199_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3570_ _3572_/A _3575_/B _3569_/X vssd1 vssd1 vccd1 vccd1 _3571_/B sky130_fd_sc_hd__o21ai_1
X_2521_ _2518_/Y _3788_/A _2521_/S vssd1 vssd1 vccd1 vccd1 _2527_/B sky130_fd_sc_hd__mux2_1
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5240_ _5445_/CLK _5240_/D vssd1 vssd1 vccd1 vccd1 _5240_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5171_ _5351_/CLK _5171_/D vssd1 vssd1 vccd1 vccd1 _5171_/Q sky130_fd_sc_hd__dfxtp_2
X_4122_ _5340_/Q _5163_/Q _4126_/S vssd1 vssd1 vccd1 vccd1 _4123_/A sky130_fd_sc_hd__mux2_1
X_4053_ _4053_/A vssd1 vssd1 vccd1 vccd1 _5138_/D sky130_fd_sc_hd__clkbuf_1
Xinput3 io_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_6
X_3004_ _3005_/A _3065_/A vssd1 vssd1 vccd1 vccd1 _3004_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4955_ _5443_/Q _4954_/C _4094_/X vssd1 vssd1 vccd1 vccd1 _4955_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_52_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3906_ _5280_/Q _3699_/A _3903_/A _5012_/Q vssd1 vssd1 vccd1 vccd1 _3906_/X sky130_fd_sc_hd__a22o_1
X_4886_ _4901_/A _4886_/B vssd1 vssd1 vccd1 vccd1 _4886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3837_ _3847_/C _3837_/B vssd1 vssd1 vccd1 vccd1 _5055_/D sky130_fd_sc_hd__nor2_1
XFILLER_137_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3768_ _3823_/A _3772_/B vssd1 vssd1 vccd1 vccd1 _3768_/Y sky130_fd_sc_hd__nand2_1
X_2719_ hold88/A _5151_/Q vssd1 vssd1 vccd1 vccd1 _2720_/C sky130_fd_sc_hd__xnor2_1
X_3699_ _3699_/A vssd1 vssd1 vccd1 vccd1 _3910_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5438_ _5446_/CLK _5438_/D vssd1 vssd1 vccd1 vccd1 _5438_/Q sky130_fd_sc_hd__dfxtp_1
X_5369_ _5369_/CLK _5369_/D vssd1 vssd1 vccd1 vccd1 _5369_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _5355_/Q _5371_/D vssd1 vssd1 vccd1 vccd1 _4744_/A sky130_fd_sc_hd__and2_1
X_4671_ _5574_/A _4669_/X _4671_/S vssd1 vssd1 vccd1 vccd1 _4672_/B sky130_fd_sc_hd__mux2_1
X_3622_ _4504_/A _3641_/B vssd1 vssd1 vccd1 vccd1 _3895_/A sky130_fd_sc_hd__nand2_1
X_3553_ _3553_/A _3553_/B vssd1 vssd1 vccd1 vccd1 _3829_/C sky130_fd_sc_hd__nor2_1
X_3484_ _3465_/Y _3481_/X _3483_/X vssd1 vssd1 vccd1 vccd1 _3484_/Y sky130_fd_sc_hd__a21oi_1
X_5223_ _5328_/CLK _5223_/D vssd1 vssd1 vccd1 vccd1 _5576_/A sky130_fd_sc_hd__dfxtp_1
X_5154_ _5160_/CLK _5154_/D vssd1 vssd1 vccd1 vccd1 _5154_/Q sky130_fd_sc_hd__dfxtp_4
X_4105_ hold46/A _4107_/C _2766_/A vssd1 vssd1 vccd1 vccd1 _4106_/B sky130_fd_sc_hd__o21ai_1
XFILLER_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5085_ _5431_/CLK _5085_/D vssd1 vssd1 vccd1 vccd1 _5085_/Q sky130_fd_sc_hd__dfxtp_1
X_4036_ _4038_/A _3470_/Y _4030_/Y vssd1 vssd1 vccd1 vccd1 _4036_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_25_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4938_ _5434_/Q _2889_/B _4938_/S vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__mux2_1
X_4869_ _5410_/Q _4869_/B vssd1 vssd1 vccd1 vccd1 _4869_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_30 _4350_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2984_ _2984_/A _2984_/B vssd1 vssd1 vccd1 vccd1 _2984_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4723_ _5333_/Q _4725_/C _4710_/B vssd1 vssd1 vccd1 vccd1 _4724_/B sky130_fd_sc_hd__o21ai_1
X_4654_ _5315_/Q _4653_/X _4662_/S vssd1 vssd1 vccd1 vccd1 _4655_/B sky130_fd_sc_hd__mux2_1
X_3605_ _3733_/B _4024_/A vssd1 vssd1 vccd1 vccd1 _3729_/B sky130_fd_sc_hd__and2_1
X_4585_ _5328_/Q vssd1 vssd1 vccd1 vccd1 _4586_/A sky130_fd_sc_hd__inv_2
X_3536_ _3665_/A _3667_/A vssd1 vssd1 vccd1 vccd1 _4285_/A sky130_fd_sc_hd__nor2_2
X_3467_ _3466_/A _2835_/Y _3465_/Y _3466_/Y vssd1 vssd1 vccd1 vccd1 _3467_/X sky130_fd_sc_hd__o211a_1
X_5206_ _5445_/CLK _5206_/D vssd1 vssd1 vccd1 vccd1 _5206_/Q sky130_fd_sc_hd__dfxtp_1
X_4001__8 _4002__9/A vssd1 vssd1 vccd1 vccd1 _5115_/CLK sky130_fd_sc_hd__inv_2
X_3398_ _3398_/A _4073_/B _4073_/C vssd1 vssd1 vccd1 vccd1 _3398_/X sky130_fd_sc_hd__or3b_1
X_5137_ _5313_/CLK _5137_/D vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
X_5068_ _5077_/CLK _5068_/D vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
X_4019_ _5126_/Q input13/X _4019_/S vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold108 hold91/X vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__clkbuf_2
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__clkbuf_2
X_4370_ _4381_/A _4370_/B vssd1 vssd1 vccd1 vccd1 _4370_/X sky130_fd_sc_hd__or2_1
X_3321_ _3321_/A _3321_/B vssd1 vssd1 vccd1 vccd1 _3344_/A sky130_fd_sc_hd__or2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3245_/X _3251_/Y _3252_/S vssd1 vssd1 vccd1 vccd1 _3309_/A sky130_fd_sc_hd__mux2_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _3646_/A _3646_/B vssd1 vssd1 vccd1 vccd1 _3183_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5435_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2967_ _2903_/C _2925_/X _2965_/X _2944_/X _2966_/X vssd1 vssd1 vccd1 vccd1 _5374_/D
+ sky130_fd_sc_hd__o221a_1
X_2898_ _2906_/A _2906_/B _2906_/C _2906_/D vssd1 vssd1 vccd1 vccd1 _2953_/C sky130_fd_sc_hd__nor4_2
X_4706_ _4714_/B vssd1 vssd1 vccd1 vccd1 _4707_/A sky130_fd_sc_hd__inv_2
X_4637_ _4655_/A _4637_/B vssd1 vssd1 vccd1 vccd1 _4638_/A sky130_fd_sc_hd__and2_1
X_4568_ _5294_/Q _4577_/B vssd1 vssd1 vccd1 vccd1 _4568_/X sky130_fd_sc_hd__or2_1
XFILLER_1_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3519_ _5207_/Q _3665_/A _3533_/A vssd1 vssd1 vccd1 vccd1 _3519_/X sky130_fd_sc_hd__o21a_1
X_4499_ _5269_/Q _5107_/Q _4519_/S vssd1 vssd1 vccd1 vccd1 _4500_/A sky130_fd_sc_hd__mux2_1
X_5488__78 vssd1 vssd1 vccd1 vccd1 _5488__78/HI _5566_/A sky130_fd_sc_hd__conb_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3870_ _3870_/A vssd1 vssd1 vccd1 vccd1 _5068_/D sky130_fd_sc_hd__clkbuf_1
X_2821_ _5131_/Q vssd1 vssd1 vccd1 vccd1 _2838_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5540_ _5540_/A _2689_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[6] sky130_fd_sc_hd__ebufn_8
X_2752_ _5112_/Q _2752_/B _2752_/C vssd1 vssd1 vccd1 vccd1 _2753_/B sky130_fd_sc_hd__or3_1
XFILLER_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2683_ _2683_/A vssd1 vssd1 vccd1 vccd1 _2683_/Y sky130_fd_sc_hd__inv_2
X_4422_ _4422_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _4422_/X sky130_fd_sc_hd__or2_1
X_4353_ _4353_/A _5252_/Q _4353_/C vssd1 vssd1 vccd1 vccd1 _4353_/X sky130_fd_sc_hd__and3_1
X_3304_ _3314_/A _3314_/B vssd1 vssd1 vccd1 vccd1 _3388_/A sky130_fd_sc_hd__xor2_2
X_4284_ _4284_/A vssd1 vssd1 vccd1 vccd1 _5212_/D sky130_fd_sc_hd__clkbuf_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _4988_/Q _4987_/Q vssd1 vssd1 vccd1 vccd1 _3559_/B sky130_fd_sc_hd__or2_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _3166_/A _3166_/B _3166_/C vssd1 vssd1 vccd1 vccd1 _3166_/Y sky130_fd_sc_hd__nand3_1
X_3097_ _3097_/A _3097_/B _3097_/C vssd1 vssd1 vccd1 vccd1 _3115_/B sky130_fd_sc_hd__or3_1
XFILLER_39_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_1_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3020_ _3020_/A _3020_/B vssd1 vssd1 vccd1 vccd1 _3021_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4971_ _2965_/X _4965_/Y _4970_/X _4902_/X vssd1 vssd1 vccd1 vccd1 _5449_/D sky130_fd_sc_hd__o211a_1
X_3922_ _5082_/Q _3909_/X _3921_/X vssd1 vssd1 vccd1 vccd1 _5082_/D sky130_fd_sc_hd__o21a_1
X_3853_ _3853_/A _3853_/B vssd1 vssd1 vccd1 vccd1 _3854_/B sky130_fd_sc_hd__xnor2_1
X_2804_ _2875_/S _2840_/A vssd1 vssd1 vccd1 vccd1 _2813_/B sky130_fd_sc_hd__nor2_1
XFILLER_32_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3784_ _5035_/Q _3767_/X _3606_/X _3784_/B2 vssd1 vssd1 vccd1 vccd1 _5035_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2735_ _5112_/Q vssd1 vssd1 vccd1 vccd1 _2739_/A sky130_fd_sc_hd__inv_2
X_2666_ _2666_/A vssd1 vssd1 vccd1 vccd1 _2671_/A sky130_fd_sc_hd__buf_2
X_5454_ _5403_/Q _5454_/D vssd1 vssd1 vccd1 vccd1 _5454_/Q sky130_fd_sc_hd__dfxtp_1
X_5385_ _5403_/Q _5385_/D vssd1 vssd1 vccd1 vccd1 _5385_/Q sky130_fd_sc_hd__dfxtp_1
X_4405_ _5201_/Q _5171_/Q _4418_/S vssd1 vssd1 vccd1 vccd1 _4406_/B sky130_fd_sc_hd__mux2_1
X_2597_ _2597_/A vssd1 vssd1 vccd1 vccd1 _2597_/Y sky130_fd_sc_hd__inv_2
X_4336_ _5576_/A _4327_/X _4348_/A vssd1 vssd1 vccd1 vccd1 _4336_/Y sky130_fd_sc_hd__a21oi_1
X_4267_ _4267_/A vssd1 vssd1 vccd1 vccd1 _5208_/D sky130_fd_sc_hd__clkbuf_1
X_5458__48 vssd1 vssd1 vccd1 vccd1 _5458__48/HI _5535_/A sky130_fd_sc_hd__conb_1
X_3218_ _3244_/C vssd1 vssd1 vccd1 vccd1 _3277_/B sky130_fd_sc_hd__buf_2
X_4198_ _4198_/A vssd1 vssd1 vccd1 vccd1 _5188_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3149_ _3166_/A _3149_/B vssd1 vssd1 vccd1 vccd1 _3150_/C sky130_fd_sc_hd__nand2_1
XFILLER_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5472__62 vssd1 vssd1 vccd1 vccd1 _5472__62/HI _5549_/A sky130_fd_sc_hd__conb_1
XFILLER_14_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2520_ _5039_/Q _5037_/Q _5036_/Q _5038_/Q vssd1 vssd1 vccd1 vccd1 _2521_/S sky130_fd_sc_hd__or4_1
X_5170_ _5351_/CLK _5170_/D vssd1 vssd1 vccd1 vccd1 _5170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4121_ _4121_/A vssd1 vssd1 vccd1 vccd1 _5162_/D sky130_fd_sc_hd__clkbuf_1
X_4052_ _2903_/B hold49/A _4054_/S vssd1 vssd1 vccd1 vccd1 _4053_/A sky130_fd_sc_hd__mux2_1
Xinput4 io_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_6
X_3003_ _3013_/B _3003_/B vssd1 vssd1 vccd1 vccd1 _3065_/A sky130_fd_sc_hd__and2_1
X_4954_ _4954_/A _4954_/B _4954_/C vssd1 vssd1 vccd1 vccd1 _5442_/D sky130_fd_sc_hd__nor3_1
XFILLER_51_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3905_ _5079_/Q _3697_/X _3700_/X _5279_/Q _3904_/X vssd1 vssd1 vccd1 vccd1 _5079_/D
+ sky130_fd_sc_hd__a221o_1
X_4885_ _5414_/Q _4888_/C vssd1 vssd1 vccd1 vccd1 _4886_/B sky130_fd_sc_hd__xnor2_1
X_3836_ _3835_/A _3834_/A _3826_/X vssd1 vssd1 vccd1 vccd1 _3837_/B sky130_fd_sc_hd__o21ai_1
X_3767_ _3767_/A vssd1 vssd1 vccd1 vccd1 _3767_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2718_ hold94/A _5152_/Q vssd1 vssd1 vccd1 vccd1 _2778_/A sky130_fd_sc_hd__xnor2_1
X_3698_ _3698_/A vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__buf_2
X_2649_ _2653_/A vssd1 vssd1 vccd1 vccd1 _2649_/Y sky130_fd_sc_hd__inv_2
X_5437_ _5437_/CLK _5437_/D vssd1 vssd1 vccd1 vccd1 _5437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5368_ _5369_/CLK _5368_/D vssd1 vssd1 vccd1 vccd1 _5368_/Q sky130_fd_sc_hd__dfxtp_1
X_5299_ _5437_/CLK _5299_/D vssd1 vssd1 vccd1 vccd1 _5299_/Q sky130_fd_sc_hd__dfxtp_1
X_4319_ _4319_/A vssd1 vssd1 vccd1 vccd1 _5220_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4670_ _4587_/A _3641_/B _4597_/Y vssd1 vssd1 vccd1 vccd1 _4671_/S sky130_fd_sc_hd__o21ba_1
X_3621_ _4328_/A _5321_/Q vssd1 vssd1 vccd1 vccd1 _3641_/B sky130_fd_sc_hd__and2_1
X_3552_ _4073_/B _4994_/Q _3559_/B _4075_/C vssd1 vssd1 vccd1 vccd1 _3553_/B sky130_fd_sc_hd__or4_1
XFILLER_6_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3483_ _3465_/A _3470_/B _3482_/X _4038_/B vssd1 vssd1 vccd1 vccd1 _3483_/X sky130_fd_sc_hd__a31o_1
X_5222_ _5369_/CLK _5222_/D vssd1 vssd1 vccd1 vccd1 _5222_/Q sky130_fd_sc_hd__dfxtp_1
X_5153_ _5328_/CLK _5153_/D vssd1 vssd1 vccd1 vccd1 _5153_/Q sky130_fd_sc_hd__dfxtp_4
X_4104_ hold46/A _4107_/C vssd1 vssd1 vccd1 vccd1 _4106_/A sky130_fd_sc_hd__and2_1
XFILLER_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5084_ _5431_/CLK _5084_/D vssd1 vssd1 vccd1 vccd1 _5084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4035_ _2822_/B _4034_/Y _4038_/A vssd1 vssd1 vccd1 vccd1 _4035_/X sky130_fd_sc_hd__a21o_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ _4937_/A vssd1 vssd1 vccd1 vccd1 _5433_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_40_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 _5641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_20 _3760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4868_ _5410_/Q _4869_/B vssd1 vssd1 vccd1 vccd1 _4875_/C sky130_fd_sc_hd__and2_1
XFILLER_20_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3819_ _5050_/Q _5049_/Q _3813_/B _5051_/Q vssd1 vssd1 vccd1 vccd1 _3820_/C sky130_fd_sc_hd__a31o_1
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4799_ _2990_/X _5390_/Q _4801_/S vssd1 vssd1 vccd1 vccd1 _4800_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2983_ _2984_/A _2984_/B vssd1 vssd1 vccd1 vccd1 _2985_/A sky130_fd_sc_hd__nor2_1
X_4722_ _5332_/Q _5333_/Q _4722_/C vssd1 vssd1 vccd1 vccd1 _4724_/A sky130_fd_sc_hd__and3_1
X_4653_ _5297_/Q _5267_/Q _4661_/S vssd1 vssd1 vccd1 vccd1 _4653_/X sky130_fd_sc_hd__mux2_1
Xinput40 la1_data_in[3] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_2
X_4584_ _5420_/Q _3075_/B _4583_/B _4583_/Y vssd1 vssd1 vccd1 vccd1 _5301_/D sky130_fd_sc_hd__a31o_1
X_3604_ _4508_/A _3604_/B vssd1 vssd1 vccd1 vccd1 _4024_/A sky130_fd_sc_hd__nor2_2
X_3535_ _3535_/A vssd1 vssd1 vccd1 vccd1 _3535_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3466_ _3466_/A _3466_/B vssd1 vssd1 vccd1 vccd1 _3466_/Y sky130_fd_sc_hd__nand2_1
X_5205_ _5445_/CLK _5205_/D vssd1 vssd1 vccd1 vccd1 _5205_/Q sky130_fd_sc_hd__dfxtp_1
X_3397_ _4994_/Q vssd1 vssd1 vccd1 vccd1 _4073_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5136_ _5313_/CLK _5136_/D vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5067_ _5077_/CLK _5067_/D vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4018_ _4018_/A vssd1 vssd1 vccd1 vccd1 _5125_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_13_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold109 hold90/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3320_ _3319_/A _3319_/B _3319_/C vssd1 vssd1 vccd1 vccd1 _3321_/B sky130_fd_sc_hd__a21oi_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3251_/A _3251_/B vssd1 vssd1 vccd1 vccd1 _3251_/Y sky130_fd_sc_hd__xnor2_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _3181_/A _3181_/B _3181_/C vssd1 vssd1 vccd1 vccd1 _3646_/C sky130_fd_sc_hd__a21oi_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2966_ _2991_/A _5230_/Q vssd1 vssd1 vccd1 vccd1 _2966_/X sky130_fd_sc_hd__or2_1
X_2897_ _5375_/Q _5374_/Q _5373_/Q vssd1 vssd1 vccd1 vccd1 _2906_/D sky130_fd_sc_hd__or3_1
X_4705_ _5330_/Q vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4636_ _5311_/Q _4635_/X _4640_/S vssd1 vssd1 vccd1 vccd1 _4637_/B sky130_fd_sc_hd__mux2_1
X_4567_ _4581_/B vssd1 vssd1 vccd1 vccd1 _4577_/B sky130_fd_sc_hd__clkbuf_1
X_3518_ _3662_/C _4363_/B vssd1 vssd1 vccd1 vccd1 _3533_/A sky130_fd_sc_hd__nand2_1
X_4498_ _4498_/A vssd1 vssd1 vccd1 vccd1 _5268_/D sky130_fd_sc_hd__clkbuf_1
X_3449_ _2866_/X _2869_/X _2838_/X vssd1 vssd1 vccd1 vccd1 _3449_/Y sky130_fd_sc_hd__a21oi_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5119_ _5119_/CLK _5119_/D vssd1 vssd1 vccd1 vccd1 _5587_/A sky130_fd_sc_hd__dfxtp_4
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5523__113 vssd1 vssd1 vccd1 vccd1 _5523__113/HI _5639_/A sky130_fd_sc_hd__conb_1
XFILLER_48_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2820_ _2827_/C vssd1 vssd1 vccd1 vccd1 _3462_/B sky130_fd_sc_hd__clkbuf_2
X_2751_ _2728_/X _2732_/X _2745_/X _2750_/X vssd1 vssd1 vccd1 vccd1 _5038_/D sky130_fd_sc_hd__o31a_1
X_2682_ _2683_/A vssd1 vssd1 vccd1 vccd1 _2682_/Y sky130_fd_sc_hd__inv_2
X_4421_ _5206_/Q _5176_/Q _4421_/S vssd1 vssd1 vccd1 vccd1 _4422_/B sky130_fd_sc_hd__mux2_1
X_4352_ _5251_/Q _5250_/Q _5249_/Q vssd1 vssd1 vccd1 vccd1 _4353_/C sky130_fd_sc_hd__nor3_1
X_3303_ _3306_/A _3408_/A _3298_/A vssd1 vssd1 vccd1 vccd1 _3314_/B sky130_fd_sc_hd__a21o_1
X_4283_ _4282_/X _5212_/Q _4288_/S vssd1 vssd1 vccd1 vccd1 _4284_/A sky130_fd_sc_hd__mux2_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _4990_/Q _3328_/A vssd1 vssd1 vccd1 vccd1 _3336_/A sky130_fd_sc_hd__nand2_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _3166_/A _3166_/B _3166_/C vssd1 vssd1 vccd1 vccd1 _3181_/B sky130_fd_sc_hd__a21o_1
XFILLER_27_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3096_ _3142_/A _3096_/B vssd1 vssd1 vccd1 vccd1 _3097_/C sky130_fd_sc_hd__xnor2_1
XFILLER_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2949_ _2913_/A _2913_/B _2938_/B _2948_/X vssd1 vssd1 vccd1 vccd1 _2961_/A sky130_fd_sc_hd__a31o_1
XFILLER_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5599_ _5599_/A _2631_/Y vssd1 vssd1 vccd1 vccd1 io_out[33] sky130_fd_sc_hd__ebufn_8
X_4619_ _4619_/A vssd1 vssd1 vccd1 vccd1 _5307_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_1_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5446_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_49_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4970_ _4965_/A _4965_/B _5602_/A vssd1 vssd1 vccd1 vccd1 _4970_/X sky130_fd_sc_hd__a21o_1
X_3921_ _5078_/Q _3904_/C _3920_/X _3911_/X vssd1 vssd1 vccd1 vccd1 _3921_/X sky130_fd_sc_hd__a211o_1
X_3852_ _3851_/A _3851_/B _3853_/B _3826_/X vssd1 vssd1 vccd1 vccd1 _5060_/D sky130_fd_sc_hd__o211a_1
X_2803_ _2795_/X _3476_/A _2816_/B vssd1 vssd1 vccd1 vccd1 _2843_/S sky130_fd_sc_hd__a21oi_2
XFILLER_32_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3783_ _5034_/Q _3767_/X _3606_/X _3783_/B2 vssd1 vssd1 vccd1 vccd1 _5034_/D sky130_fd_sc_hd__a22o_1
XFILLER_9_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2734_ _2734_/A _5114_/Q vssd1 vssd1 vccd1 vccd1 _2737_/C sky130_fd_sc_hd__nor2_1
X_2665_ _2665_/A vssd1 vssd1 vccd1 vccd1 _2665_/Y sky130_fd_sc_hd__inv_2
X_5453_ _5403_/Q _5453_/D vssd1 vssd1 vccd1 vccd1 _5453_/Q sky130_fd_sc_hd__dfxtp_1
X_2596_ _2597_/A vssd1 vssd1 vccd1 vccd1 _2596_/Y sky130_fd_sc_hd__inv_2
X_5384_ _5403_/Q _5384_/D vssd1 vssd1 vccd1 vccd1 _5384_/Q sky130_fd_sc_hd__dfxtp_4
X_4404_ _4421_/S vssd1 vssd1 vccd1 vccd1 _4418_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_5_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4335_ _5267_/Q _3915_/X _4329_/X _4334_/X vssd1 vssd1 vccd1 vccd1 _4335_/Y sky130_fd_sc_hd__a211oi_1
X_4266_ _4265_/X _5208_/Q _4266_/S vssd1 vssd1 vccd1 vccd1 _4267_/A sky130_fd_sc_hd__mux2_1
X_3217_ _5052_/Q vssd1 vssd1 vccd1 vccd1 _3829_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4197_ _4196_/X _5188_/Q _4197_/S vssd1 vssd1 vccd1 vccd1 _4198_/A sky130_fd_sc_hd__mux2_1
X_3148_ _3148_/A _3148_/B vssd1 vssd1 vccd1 vccd1 _3149_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3079_ _3142_/A _3079_/B vssd1 vssd1 vccd1 vccd1 _3083_/B sky130_fd_sc_hd__xnor2_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4120_ _5339_/Q _5162_/Q _4126_/S vssd1 vssd1 vccd1 vccd1 _4121_/A sky130_fd_sc_hd__mux2_1
X_4051_ _4051_/A vssd1 vssd1 vccd1 vccd1 _5137_/D sky130_fd_sc_hd__clkbuf_1
Xinput5 io_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_6
X_3002_ _3002_/A _3002_/B vssd1 vssd1 vccd1 vccd1 _3003_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4953_ _5442_/Q _4953_/B _4953_/C vssd1 vssd1 vccd1 vccd1 _4954_/C sky130_fd_sc_hd__and3_1
XFILLER_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3904_ _5013_/Q _3959_/S _3904_/C vssd1 vssd1 vccd1 vccd1 _3904_/X sky130_fd_sc_hd__and3_1
X_4884_ _4884_/A vssd1 vssd1 vccd1 vccd1 _4884_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3835_ _3835_/A _3835_/B _3835_/C vssd1 vssd1 vccd1 vccd1 _3847_/C sky130_fd_sc_hd__and3_1
X_3766_ _5028_/Q _3602_/X _3740_/X _3765_/X vssd1 vssd1 vccd1 vccd1 _5028_/D sky130_fd_sc_hd__a22o_1
X_2717_ hold46/A _5153_/Q vssd1 vssd1 vccd1 vccd1 _2717_/X sky130_fd_sc_hd__xor2_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3697_ _3697_/A vssd1 vssd1 vccd1 vccd1 _3697_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5436_ _5436_/CLK _5436_/D vssd1 vssd1 vccd1 vccd1 _5436_/Q sky130_fd_sc_hd__dfxtp_1
X_2648_ _2666_/A vssd1 vssd1 vccd1 vccd1 _2653_/A sky130_fd_sc_hd__buf_2
X_2579_ input1/X vssd1 vssd1 vccd1 vccd1 _2604_/A sky130_fd_sc_hd__buf_4
X_5367_ _5369_/CLK _5367_/D vssd1 vssd1 vccd1 vccd1 _5367_/Q sky130_fd_sc_hd__dfxtp_1
X_5298_ _5437_/CLK _5298_/D vssd1 vssd1 vccd1 vccd1 _5298_/Q sky130_fd_sc_hd__dfxtp_1
X_4318_ _4317_/X _5220_/Q _4324_/S vssd1 vssd1 vccd1 vccd1 _4319_/A sky130_fd_sc_hd__mux2_1
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4249_ _4252_/A _4249_/B vssd1 vssd1 vccd1 vccd1 _4250_/A sky130_fd_sc_hd__and2_1
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3620_ _5322_/Q vssd1 vssd1 vccd1 vccd1 _4328_/A sky130_fd_sc_hd__inv_2
X_3551_ _3563_/A _3551_/B _3551_/C _3572_/B vssd1 vssd1 vccd1 vccd1 _4075_/C sky130_fd_sc_hd__or4b_1
XFILLER_6_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3482_ _5019_/Q _5022_/Q _5021_/Q _5020_/Q _2833_/A _2846_/A vssd1 vssd1 vccd1 vccd1
+ _3482_/X sky130_fd_sc_hd__mux4_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5221_ _5369_/CLK _5221_/D vssd1 vssd1 vccd1 vccd1 _5221_/Q sky130_fd_sc_hd__dfxtp_1
X_5152_ _5328_/CLK _5152_/D vssd1 vssd1 vccd1 vccd1 _5152_/Q sky130_fd_sc_hd__dfxtp_4
X_4103_ _4107_/C _4103_/B vssd1 vssd1 vccd1 vccd1 _5157_/D sky130_fd_sc_hd__nor2_1
X_5083_ _5431_/CLK _5083_/D vssd1 vssd1 vccd1 vccd1 _5083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4034_ _4034_/A _4034_/B vssd1 vssd1 vccd1 vccd1 _4034_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4936_ _5433_/Q _5384_/Q _4938_/S vssd1 vssd1 vccd1 vccd1 _4937_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_32 _5641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 _3760_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4867_ _5377_/D _4863_/X _4866_/Y _4861_/X vssd1 vssd1 vccd1 vccd1 _5409_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_10 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ _5050_/Q _5051_/Q _3818_/C vssd1 vssd1 vccd1 vccd1 _3820_/B sky130_fd_sc_hd__nand3_1
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4798_ _4798_/A vssd1 vssd1 vccd1 vccd1 _5389_/D sky130_fd_sc_hd__clkbuf_1
X_3749_ _3772_/B _3749_/B vssd1 vssd1 vccd1 vccd1 _3749_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5419_ _5445_/CLK _5419_/D vssd1 vssd1 vccd1 vccd1 _5419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2982_ _3130_/A _2982_/B vssd1 vssd1 vccd1 vccd1 _2984_/B sky130_fd_sc_hd__xnor2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _4721_/A vssd1 vssd1 vccd1 vccd1 _5332_/D sky130_fd_sc_hd__clkbuf_1
X_4652_ _4652_/A vssd1 vssd1 vccd1 vccd1 _5314_/D sky130_fd_sc_hd__clkbuf_1
X_3603_ _3754_/A vssd1 vssd1 vccd1 vccd1 _3606_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput30 la1_data_in[1] vssd1 vssd1 vccd1 vccd1 _2907_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput41 la1_data_in[4] vssd1 vssd1 vccd1 vccd1 _2977_/B sky130_fd_sc_hd__clkbuf_2
X_4583_ _4583_/A _4583_/B vssd1 vssd1 vccd1 vccd1 _4583_/Y sky130_fd_sc_hd__nor2_1
X_3534_ _3658_/B _3534_/B vssd1 vssd1 vccd1 vccd1 _3535_/A sky130_fd_sc_hd__or2_1
X_3465_ _3465_/A _3470_/B vssd1 vssd1 vccd1 vccd1 _3465_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5204_ _5245_/CLK _5204_/D vssd1 vssd1 vccd1 vccd1 _5204_/Q sky130_fd_sc_hd__dfxtp_1
X_3396_ _3396_/A _3396_/B vssd1 vssd1 vccd1 vccd1 _3396_/Y sky130_fd_sc_hd__nor2_1
X_5135_ _5313_/CLK _5135_/D vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
X_5066_ _5077_/CLK _5066_/D vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
X_4017_ _5125_/Q input12/X _4019_/S vssd1 vssd1 vccd1 vccd1 _4018_/A sky130_fd_sc_hd__mux2_1
XFILLER_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xsoc.spi_video_ram_1.write_fifo.dffrf _5160_/CLK _3707_/C_N _3746_/A0 _3753_/A0 _3760_/A0
+ _3764_/A0 _3769_/A0 _3773_/A0 _3608_/B2 _3607_/B2 _3784_/B2 _3783_/B2 _3713_/C_N
+ _3782_/B2 _3779_/A2 _3776_/A2 _3773_/A1 _3769_/A1 _3764_/A1 _3760_/A1 _3753_/A1
+ _3746_/A1 soc.spi_video_ram_1.write_fifo.dffrf/DA[29] _3718_/A soc.spi_video_ram_1.write_fifo.dffrf/DA[30]
+ soc.spi_video_ram_1.write_fifo.dffrf/DA[31] _3722_/A _3724_/A _3726_/C_N _3728_/A1
+ _3734_/A _3737_/A1 _3742_/A1 soc.spi_video_ram_1.write_fifo.dffrf/DB[0] soc.spi_video_ram_1.write_fifo.dffrf/DB[10]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[11] soc.spi_video_ram_1.write_fifo.dffrf/DB[12]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[13] soc.spi_video_ram_1.write_fifo.dffrf/DB[14]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[15] soc.spi_video_ram_1.write_fifo.dffrf/DB[16]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[17] soc.spi_video_ram_1.write_fifo.dffrf/DB[18]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[19] soc.spi_video_ram_1.write_fifo.dffrf/DB[1]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[20] soc.spi_video_ram_1.write_fifo.dffrf/DB[21]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[22] soc.spi_video_ram_1.write_fifo.dffrf/DB[23]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[24] soc.spi_video_ram_1.write_fifo.dffrf/DB[25]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[26] soc.spi_video_ram_1.write_fifo.dffrf/DB[27]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[28] soc.spi_video_ram_1.write_fifo.dffrf/DB[29]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[2] soc.spi_video_ram_1.write_fifo.dffrf/DB[30]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[31] soc.spi_video_ram_1.write_fifo.dffrf/DB[3]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[4] soc.spi_video_ram_1.write_fifo.dffrf/DB[5]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[6] soc.spi_video_ram_1.write_fifo.dffrf/DB[7]
+ soc.spi_video_ram_1.write_fifo.dffrf/DB[8] soc.spi_video_ram_1.write_fifo.dffrf/DB[9]
+ hold131/X hold9/X hold30/X hold21/X hold12/X hold6/X hold18/X hold57/X hold60/X
+ hold75/X hold51/X hold127/X hold81/X hold72/X hold54/X hold63/X hold87/X hold66/X
+ hold78/X hold69/X hold84/X _5526__116/LO hold128/X _5527__117/LO _5528__118/LO hold42/X
+ hold27/X hold36/X hold33/X hold24/X hold15/X hold3/X hold122/X hold124/X hold48/X
+ hold45/X hold39/X _5529__119/LO _5530__120/LO _5531__121/LO _5532__122/LO _5533__123/LO
+ hold114/X hold119/X hold116/X hold108/X hold136/X vssd1 vccd1 _5456__125/HI DFFRF_2R1W
XFILLER_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4919_ _5425_/Q _5376_/Q _4927_/S vssd1 vssd1 vccd1 vccd1 _4920_/A sky130_fd_sc_hd__mux2_1
XFILLER_21_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5502__92 vssd1 vssd1 vccd1 vccd1 _5502__92/HI _5605_/A sky130_fd_sc_hd__conb_1
XFILLER_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _3250_/A _3249_/X vssd1 vssd1 vccd1 vccd1 _3251_/B sky130_fd_sc_hd__or2b_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _3181_/A _3181_/B _3181_/C vssd1 vssd1 vccd1 vccd1 _3181_/X sky130_fd_sc_hd__and3_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4704_ _5329_/Q vssd1 vssd1 vccd1 vccd1 _4714_/A sky130_fd_sc_hd__clkbuf_1
X_2965_ _4831_/C vssd1 vssd1 vccd1 vccd1 _2965_/X sky130_fd_sc_hd__clkbuf_4
X_2896_ _5381_/Q _5380_/Q _5386_/Q _5385_/Q vssd1 vssd1 vccd1 vccd1 _2906_/C sky130_fd_sc_hd__or4bb_2
XFILLER_30_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4635_ _5293_/Q _5263_/Q _4639_/S vssd1 vssd1 vccd1 vccd1 _4635_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5444_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4566_ _4566_/A vssd1 vssd1 vccd1 vccd1 _4566_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3517_ _4730_/A _5247_/Q vssd1 vssd1 vccd1 vccd1 _4363_/B sky130_fd_sc_hd__nor2_2
X_4497_ _5268_/Q _5106_/Q _4519_/S vssd1 vssd1 vccd1 vccd1 _4498_/A sky130_fd_sc_hd__mux2_1
X_3448_ _4034_/B _3476_/B vssd1 vssd1 vccd1 vccd1 _3448_/Y sky130_fd_sc_hd__xnor2_2
X_3379_ _3379_/A _3379_/B vssd1 vssd1 vccd1 vccd1 _3380_/B sky130_fd_sc_hd__nor2_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5118_/CLK _5118_/D vssd1 vssd1 vccd1 vccd1 _5118_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5049_ _5051_/CLK _5049_/D vssd1 vssd1 vccd1 vccd1 _5049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5479__69 vssd1 vssd1 vccd1 vccd1 _5479__69/HI _5556_/A sky130_fd_sc_hd__conb_1
XFILLER_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2750_ _4571_/A vssd1 vssd1 vccd1 vccd1 _2750_/X sky130_fd_sc_hd__buf_2
X_2681_ _2683_/A vssd1 vssd1 vccd1 vccd1 _2681_/Y sky130_fd_sc_hd__inv_2
X_4420_ _5242_/Q _4402_/X _4419_/X _4416_/X vssd1 vssd1 vccd1 vccd1 _5242_/D sky130_fd_sc_hd__o211a_1
X_4351_ _5253_/Q vssd1 vssd1 vccd1 vccd1 _4353_/A sky130_fd_sc_hd__inv_2
X_3302_ _3302_/A _4074_/B vssd1 vssd1 vccd1 vccd1 _3408_/A sky130_fd_sc_hd__nand2_1
X_4282_ _5208_/Q _4275_/X _4281_/X vssd1 vssd1 vccd1 vccd1 _4282_/X sky130_fd_sc_hd__a21o_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3233_ _3238_/A _3233_/B vssd1 vssd1 vccd1 vccd1 _3268_/A sky130_fd_sc_hd__xnor2_2
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _3181_/A _3164_/B vssd1 vssd1 vccd1 vccd1 _3166_/C sky130_fd_sc_hd__nand2_1
X_5493__83 vssd1 vssd1 vccd1 vccd1 _5493__83/HI _5571_/A sky130_fd_sc_hd__conb_1
X_3095_ _3176_/A _3095_/B vssd1 vssd1 vccd1 vccd1 _3096_/B sky130_fd_sc_hd__and2_1
XFILLER_35_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2948_ _2948_/A _2948_/B _2948_/C vssd1 vssd1 vccd1 vccd1 _2948_/X sky130_fd_sc_hd__and3_1
XFILLER_13_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4618_ _4632_/A _4618_/B vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__and2_1
X_2879_ _2854_/Y _2838_/X _2862_/X _2878_/X vssd1 vssd1 vccd1 vccd1 _3489_/B sky130_fd_sc_hd__a31o_1
X_5598_ _5598_/A _2630_/Y vssd1 vssd1 vccd1 vccd1 io_out[32] sky130_fd_sc_hd__ebufn_8
X_4549_ _5288_/Q _5435_/Q _4549_/S vssd1 vssd1 vccd1 vccd1 _4550_/A sky130_fd_sc_hd__mux2_1
XFILLER_1_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3920_ _5256_/Q _3919_/X _3910_/A _5282_/Q vssd1 vssd1 vccd1 vccd1 _3920_/X sky130_fd_sc_hd__a22o_1
XFILLER_44_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3851_ _3851_/A _3851_/B vssd1 vssd1 vccd1 vccd1 _3853_/B sky130_fd_sc_hd__nand2_1
X_3782_ _5033_/Q _3767_/X _3606_/X _3782_/B2 vssd1 vssd1 vccd1 vccd1 _5033_/D sky130_fd_sc_hd__a22o_1
X_2802_ _2870_/B _2824_/S vssd1 vssd1 vccd1 vccd1 _2816_/B sky130_fd_sc_hd__nor2_1
X_2733_ _5040_/Q vssd1 vssd1 vccd1 vccd1 _3750_/A sky130_fd_sc_hd__buf_2
X_2664_ _2665_/A vssd1 vssd1 vccd1 vccd1 _2664_/Y sky130_fd_sc_hd__inv_2
X_5452_ _5403_/Q _5452_/D vssd1 vssd1 vccd1 vccd1 _5452_/Q sky130_fd_sc_hd__dfxtp_1
X_2595_ _2597_/A vssd1 vssd1 vccd1 vccd1 _2595_/Y sky130_fd_sc_hd__inv_2
X_5383_ _5403_/Q _5383_/D vssd1 vssd1 vccd1 vccd1 _5383_/Q sky130_fd_sc_hd__dfxtp_4
X_4403_ _4422_/A vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__clkbuf_1
X_4334_ _4693_/B _4330_/X _4333_/X _3942_/B _5089_/Q vssd1 vssd1 vccd1 vccd1 _4334_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4265_ _5184_/Q _3682_/D _4264_/X _5010_/Q vssd1 vssd1 vccd1 vccd1 _4265_/X sky130_fd_sc_hd__a22o_1
X_3216_ _3216_/A _3244_/C _5440_/Q vssd1 vssd1 vccd1 vccd1 _3221_/A sky130_fd_sc_hd__or3b_1
X_4196_ _5412_/Q _5363_/Q _4199_/S vssd1 vssd1 vccd1 vccd1 _4196_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3147_ _3099_/A _3115_/X _3144_/X _3146_/X _3132_/X vssd1 vssd1 vccd1 vccd1 _3150_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_27_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3078_ _3176_/A _3078_/B vssd1 vssd1 vccd1 vccd1 _3079_/B sky130_fd_sc_hd__and2_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _2903_/C hold73/A _4054_/S vssd1 vssd1 vccd1 vccd1 _4051_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput6 io_in[16] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_6
XFILLER_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3001_ _2984_/Y _2987_/B _2985_/A vssd1 vssd1 vccd1 vccd1 _3005_/A sky130_fd_sc_hd__a21o_1
XFILLER_52_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5463__53 vssd1 vssd1 vccd1 vccd1 _5463__53/HI _5540_/A sky130_fd_sc_hd__conb_1
XFILLER_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4952_ _4953_/B _4953_/C _5442_/Q vssd1 vssd1 vccd1 vccd1 _4954_/B sky130_fd_sc_hd__a21oi_1
XFILLER_51_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4883_ _5381_/D _4863_/X _4881_/Y _4882_/X vssd1 vssd1 vccd1 vccd1 _5413_/D sky130_fd_sc_hd__o211a_1
X_3903_ _3903_/A vssd1 vssd1 vccd1 vccd1 _3904_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3834_ _3834_/A _3834_/B vssd1 vssd1 vccd1 vccd1 _5054_/D sky130_fd_sc_hd__nor2_1
X_3765_ _3741_/X _3277_/Y _3764_/X _3606_/A vssd1 vssd1 vccd1 vccd1 _3765_/X sky130_fd_sc_hd__a22o_1
X_2716_ hold43/A _5154_/Q vssd1 vssd1 vccd1 vccd1 _2780_/A sky130_fd_sc_hd__xnor2_1
X_3696_ _3911_/A vssd1 vssd1 vccd1 vccd1 _3697_/A sky130_fd_sc_hd__clkbuf_2
X_5435_ _5435_/CLK _5435_/D vssd1 vssd1 vccd1 vccd1 _5435_/Q sky130_fd_sc_hd__dfxtp_1
X_2647_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2647_/Y sky130_fd_sc_hd__inv_2
X_2578_ _2578_/A vssd1 vssd1 vccd1 vccd1 _2578_/Y sky130_fd_sc_hd__inv_2
X_5366_ _5371_/CLK _5366_/D vssd1 vssd1 vccd1 vccd1 _5366_/Q sky130_fd_sc_hd__dfxtp_1
X_5297_ _5328_/CLK _5297_/D vssd1 vssd1 vccd1 vccd1 _5297_/Q sky130_fd_sc_hd__dfxtp_1
X_4317_ _5170_/Q _3537_/X _3674_/B _4316_/X vssd1 vssd1 vccd1 vccd1 _4317_/X sky130_fd_sc_hd__a211o_1
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4248_ _5203_/Q _5199_/Q _4251_/S vssd1 vssd1 vccd1 vccd1 _4249_/B sky130_fd_sc_hd__mux2_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4179_ _5407_/Q _5358_/Q _4182_/S vssd1 vssd1 vccd1 vccd1 _4179_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3550_ _5585_/A _3677_/B _3549_/X _2761_/X vssd1 vssd1 vccd1 vccd1 _4986_/D sky130_fd_sc_hd__a211o_1
X_3481_ _3480_/X _5018_/Q _5017_/Q _5016_/Q _2795_/X _2846_/A vssd1 vssd1 vccd1 vccd1
+ _3481_/X sky130_fd_sc_hd__mux4_1
XFILLER_6_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5220_ _5245_/CLK _5220_/D vssd1 vssd1 vccd1 vccd1 _5220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5151_ _5328_/CLK _5151_/D vssd1 vssd1 vccd1 vccd1 _5151_/Q sky130_fd_sc_hd__dfxtp_4
X_4102_ hold94/A _4100_/A _4081_/X vssd1 vssd1 vccd1 vccd1 _4103_/B sky130_fd_sc_hd__o21ai_1
X_5082_ _5431_/CLK _5082_/D vssd1 vssd1 vccd1 vccd1 _5082_/Q sky130_fd_sc_hd__dfxtp_1
X_4033_ _4033_/A _4033_/B vssd1 vssd1 vccd1 vccd1 _5129_/D sky130_fd_sc_hd__nand2_1
XFILLER_37_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4935_ _4935_/A vssd1 vssd1 vccd1 vccd1 _5432_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_22 _3753_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4866_ _4869_/B _4865_/Y _4851_/X vssd1 vssd1 vccd1 vccd1 _4866_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_11 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_33 _4508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3817_ _5050_/Q _3818_/C _3816_/Y vssd1 vssd1 vccd1 vccd1 _5050_/D sky130_fd_sc_hd__a21oi_1
X_4797_ _2965_/X _5389_/Q _4801_/S vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__mux2_1
X_3748_ _5025_/Q _3602_/X _3740_/X _3747_/X vssd1 vssd1 vccd1 vccd1 _5025_/D sky130_fd_sc_hd__a22o_1
XFILLER_21_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3679_ _4324_/S vssd1 vssd1 vccd1 vccd1 _4266_/S sky130_fd_sc_hd__clkbuf_2
X_5418_ _5403_/Q _5418_/D vssd1 vssd1 vccd1 vccd1 _5418_/Q sky130_fd_sc_hd__dfxtp_1
X_5349_ _5353_/CLK _5349_/D vssd1 vssd1 vccd1 vccd1 _5349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_137_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2981_ _3155_/B _2903_/B _2976_/X _2979_/X _3129_/A vssd1 vssd1 vccd1 vccd1 _2982_/B
+ sky130_fd_sc_hd__o221a_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4720_ _4725_/C _4720_/B _4720_/C vssd1 vssd1 vccd1 vccd1 _4721_/A sky130_fd_sc_hd__and3b_1
X_4651_ _4655_/A _4651_/B vssd1 vssd1 vccd1 vccd1 _4652_/A sky130_fd_sc_hd__and2_1
X_3602_ _3767_/A vssd1 vssd1 vccd1 vccd1 _3602_/X sky130_fd_sc_hd__clkbuf_2
Xinput31 la1_data_in[20] vssd1 vssd1 vccd1 vccd1 _5347_/D sky130_fd_sc_hd__clkbuf_1
Xinput20 la1_data_in[10] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__clkbuf_1
XFILLER_30_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput42 la1_data_in[5] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_2
X_4582_ _5296_/Q _4566_/A _4581_/X _4350_/X vssd1 vssd1 vccd1 vccd1 _5300_/D sky130_fd_sc_hd__o211a_1
X_3533_ _3533_/A _3533_/B vssd1 vssd1 vccd1 vccd1 _3534_/B sky130_fd_sc_hd__nand2_1
X_3464_ _3464_/A _3464_/B vssd1 vssd1 vccd1 vccd1 _3470_/B sky130_fd_sc_hd__or2_1
X_5203_ _5446_/CLK _5203_/D vssd1 vssd1 vccd1 vccd1 _5203_/Q sky130_fd_sc_hd__dfxtp_1
X_5134_ _5313_/CLK _5134_/D vssd1 vssd1 vccd1 vccd1 _5134_/Q sky130_fd_sc_hd__dfxtp_2
X_3395_ _3395_/A _3394_/X vssd1 vssd1 vccd1 vccd1 _3395_/X sky130_fd_sc_hd__or2b_1
X_5065_ _5077_/CLK _5065_/D vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfxtp_1
X_4016_ _4016_/A vssd1 vssd1 vccd1 vccd1 _5124_/D sky130_fd_sc_hd__clkbuf_1
X_3996__4 _3996__4/A vssd1 vssd1 vccd1 vccd1 _5111_/CLK sky130_fd_sc_hd__inv_2
XFILLER_12_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4918_ _4940_/S vssd1 vssd1 vccd1 vccd1 _4927_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_40_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4849_ _5404_/Q _5405_/Q _5406_/Q vssd1 vssd1 vccd1 vccd1 _4849_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_57_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _3646_/B _3180_/B vssd1 vssd1 vccd1 vccd1 _3181_/C sky130_fd_sc_hd__or2_1
XFILLER_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2964_ _3023_/A _2964_/B vssd1 vssd1 vccd1 vccd1 _4831_/C sky130_fd_sc_hd__xor2_1
X_4703_ _4586_/A _4700_/C _4702_/X _4350_/X vssd1 vssd1 vccd1 vccd1 _5328_/D sky130_fd_sc_hd__o211a_1
X_2895_ _5383_/Q _5382_/Q _5384_/Q _5377_/Q vssd1 vssd1 vccd1 vccd1 _2906_/B sky130_fd_sc_hd__or4_2
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4634_ _4634_/A vssd1 vssd1 vccd1 vccd1 _4655_/A sky130_fd_sc_hd__clkbuf_1
X_4565_ _5289_/Q _4552_/X _4564_/X _4558_/X vssd1 vssd1 vccd1 vccd1 _5293_/D sky130_fd_sc_hd__o211a_1
X_3516_ _5246_/Q _3532_/A vssd1 vssd1 vccd1 vccd1 _3665_/A sky130_fd_sc_hd__nand2_2
X_4496_ _4496_/A vssd1 vssd1 vccd1 vccd1 _5267_/D sky130_fd_sc_hd__clkbuf_1
X_3447_ _3447_/A vssd1 vssd1 vccd1 vccd1 _5593_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3378_ _3563_/B _3378_/B vssd1 vssd1 vccd1 vccd1 _3378_/Y sky130_fd_sc_hd__nor2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5117_/CLK _5117_/D vssd1 vssd1 vccd1 vccd1 _5117_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5048_ _5051_/CLK _5048_/D vssd1 vssd1 vccd1 vccd1 _5048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2680_ _2683_/A vssd1 vssd1 vccd1 vccd1 _2680_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4350_ _4350_/A vssd1 vssd1 vccd1 vccd1 _4350_/X sky130_fd_sc_hd__buf_4
X_3301_ _3396_/A _3305_/B vssd1 vssd1 vccd1 vccd1 _3306_/A sky130_fd_sc_hd__nor2_1
X_4281_ _5162_/Q _3541_/X _4276_/X _5188_/Q vssd1 vssd1 vccd1 vccd1 _4281_/X sky130_fd_sc_hd__a22o_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3252_/S _3221_/B _3231_/X vssd1 vssd1 vccd1 vccd1 _3233_/B sky130_fd_sc_hd__a21bo_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _3163_/A _3163_/B vssd1 vssd1 vccd1 vccd1 _3164_/B sky130_fd_sc_hd__nand2_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3094_ _3074_/X _5381_/Q _3076_/A _5312_/Q vssd1 vssd1 vccd1 vccd1 _3095_/B sky130_fd_sc_hd__a22o_1
XFILLER_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2947_ _2902_/X _2925_/X _2942_/X _2944_/X _2946_/X vssd1 vssd1 vccd1 vccd1 _5373_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4617_ _5307_/Q _4616_/X _4617_/S vssd1 vssd1 vccd1 vccd1 _4618_/B sky130_fd_sc_hd__mux2_1
X_2878_ _2838_/A _2878_/B vssd1 vssd1 vccd1 vccd1 _2878_/X sky130_fd_sc_hd__and2b_1
X_5597_ _5597_/A _2628_/Y vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__ebufn_8
X_4548_ _4548_/A vssd1 vssd1 vccd1 vccd1 _5287_/D sky130_fd_sc_hd__clkbuf_1
X_4479_ _5260_/Q _5098_/Q _4481_/S vssd1 vssd1 vccd1 vccd1 _4480_/A sky130_fd_sc_hd__mux2_1
XFILLER_58_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3850_ _3850_/A vssd1 vssd1 vccd1 vccd1 _5059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3781_ _3781_/A vssd1 vssd1 vccd1 vccd1 _5032_/D sky130_fd_sc_hd__clkbuf_1
X_2801_ _2875_/S _2840_/A vssd1 vssd1 vccd1 vccd1 _2824_/S sky130_fd_sc_hd__and2_1
XFILLER_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2732_ _2706_/A _2706_/B _3726_/A _3596_/A vssd1 vssd1 vccd1 vccd1 _2732_/X sky130_fd_sc_hd__o211a_1
XFILLER_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2663_ _2665_/A vssd1 vssd1 vccd1 vccd1 _2663_/Y sky130_fd_sc_hd__inv_2
X_5451_ _5403_/Q _5451_/D vssd1 vssd1 vccd1 vccd1 _5451_/Q sky130_fd_sc_hd__dfxtp_1
X_2594_ _2597_/A vssd1 vssd1 vccd1 vccd1 _2594_/Y sky130_fd_sc_hd__inv_2
X_5382_ _5403_/Q _5382_/D vssd1 vssd1 vccd1 vccd1 _5382_/Q sky130_fd_sc_hd__dfxtp_4
X_4402_ _4402_/A vssd1 vssd1 vccd1 vccd1 _4402_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4333_ _4586_/C _4333_/B _4586_/D vssd1 vssd1 vccd1 vccd1 _4333_/X sky130_fd_sc_hd__or3_1
X_4264_ _4275_/A vssd1 vssd1 vccd1 vccd1 _4264_/X sky130_fd_sc_hd__clkbuf_2
X_3215_ _3213_/Y _3260_/D _3260_/A vssd1 vssd1 vccd1 vccd1 _3215_/X sky130_fd_sc_hd__mux2_1
X_4195_ _4195_/A vssd1 vssd1 vccd1 vccd1 _5187_/D sky130_fd_sc_hd__clkbuf_1
X_3146_ _3146_/A _3146_/B vssd1 vssd1 vccd1 vccd1 _3146_/X sky130_fd_sc_hd__or2_1
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3077_ _3074_/X _5380_/Q _3076_/X _5311_/Q vssd1 vssd1 vccd1 vccd1 _3078_/B sky130_fd_sc_hd__a22o_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5513__103 vssd1 vssd1 vccd1 vccd1 _5513__103/HI _5624_/A sky130_fd_sc_hd__conb_1
XFILLER_11_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3979_ _5100_/Q _3976_/X _3973_/X _4832_/C vssd1 vssd1 vccd1 vccd1 _5100_/D sky130_fd_sc_hd__a22o_1
XFILLER_136_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput7 io_in[17] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_6
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3000_ _3002_/A _3002_/B vssd1 vssd1 vccd1 vccd1 _3013_/B sky130_fd_sc_hd__or2_1
XFILLER_37_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4951_ _4953_/B _4953_/C _4950_/Y vssd1 vssd1 vccd1 vccd1 _5441_/D sky130_fd_sc_hd__o21a_1
XFILLER_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4882_ _4902_/A vssd1 vssd1 vccd1 vccd1 _4882_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3902_ _3902_/A vssd1 vssd1 vccd1 vccd1 _5078_/D sky130_fd_sc_hd__clkbuf_1
X_3833_ _3835_/B _3835_/C _3826_/X vssd1 vssd1 vccd1 vccd1 _3834_/B sky130_fd_sc_hd__o21ai_1
XFILLER_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3764_ _3764_/A0 _3764_/A1 _3764_/S vssd1 vssd1 vccd1 vccd1 _3764_/X sky130_fd_sc_hd__mux2_1
X_2715_ hold37/A _5155_/Q vssd1 vssd1 vccd1 vccd1 _2782_/A sky130_fd_sc_hd__xnor2_1
X_3695_ _3698_/A _4347_/S vssd1 vssd1 vccd1 vccd1 _3911_/A sky130_fd_sc_hd__nand2_1
X_5434_ _5435_/CLK _5434_/D vssd1 vssd1 vccd1 vccd1 _5434_/Q sky130_fd_sc_hd__dfxtp_1
X_2646_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2646_/Y sky130_fd_sc_hd__inv_2
X_2577_ _2578_/A vssd1 vssd1 vccd1 vccd1 _2577_/Y sky130_fd_sc_hd__inv_2
X_5365_ _5444_/CLK _5365_/D vssd1 vssd1 vccd1 vccd1 _5365_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4316_ _4355_/A _3667_/A _4220_/C _3543_/B _5216_/Q vssd1 vssd1 vccd1 vccd1 _4316_/X
+ sky130_fd_sc_hd__o32a_1
X_5296_ _5437_/CLK _5296_/D vssd1 vssd1 vccd1 vccd1 _5296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4247_ _4247_/A vssd1 vssd1 vccd1 vccd1 _5202_/D sky130_fd_sc_hd__clkbuf_1
X_4178_ _4178_/A vssd1 vssd1 vccd1 vccd1 _5182_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3129_ _3129_/A _3129_/B vssd1 vssd1 vccd1 vccd1 _3130_/B sky130_fd_sc_hd__and2_1
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_0_0_wb_clk_i clkbuf_2_1_0_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5509__99 vssd1 vssd1 vccd1 vccd1 _5509__99/HI _5612_/A sky130_fd_sc_hd__conb_1
XFILLER_136_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3480_ _5015_/Q _3480_/B vssd1 vssd1 vccd1 vccd1 _3480_/X sky130_fd_sc_hd__and2_1
XFILLER_6_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5150_ _5439_/CLK _5150_/D vssd1 vssd1 vccd1 vccd1 _5150_/Q sky130_fd_sc_hd__dfxtp_1
X_4101_ hold94/A hold88/A _4101_/C vssd1 vssd1 vccd1 vccd1 _4107_/C sky130_fd_sc_hd__and3_1
X_5081_ _5431_/CLK _5081_/D vssd1 vssd1 vccd1 vccd1 _5081_/Q sky130_fd_sc_hd__dfxtp_1
X_4032_ _4034_/A _4041_/B vssd1 vssd1 vccd1 vccd1 _4033_/B sky130_fd_sc_hd__xnor2_1
XFILLER_49_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4934_ _5432_/Q _5383_/Q _4938_/S vssd1 vssd1 vccd1 vccd1 _4935_/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_19_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5126_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_23 _3753_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4865_ _5408_/Q _4864_/C _5409_/Q vssd1 vssd1 vccd1 vccd1 _4865_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_12 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3816_ _5050_/Q _3818_/C _3800_/X vssd1 vssd1 vccd1 vccd1 _3816_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4796_ _4796_/A vssd1 vssd1 vccd1 vccd1 _5388_/D sky130_fd_sc_hd__clkbuf_1
X_3747_ _3741_/X _3745_/Y _3746_/X _3606_/A vssd1 vssd1 vccd1 vccd1 _3747_/X sky130_fd_sc_hd__a22o_1
XFILLER_137_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3678_ _4292_/A vssd1 vssd1 vccd1 vccd1 _4324_/S sky130_fd_sc_hd__clkbuf_2
X_2629_ _2635_/A vssd1 vssd1 vccd1 vccd1 _2634_/A sky130_fd_sc_hd__buf_2
X_5417_ _5403_/Q _5417_/D vssd1 vssd1 vccd1 vccd1 _5417_/Q sky130_fd_sc_hd__dfxtp_1
X_5348_ _5351_/CLK _5348_/D vssd1 vssd1 vccd1 vccd1 _5348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5279_ _5430_/CLK _5279_/D vssd1 vssd1 vccd1 vccd1 _5279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2980_ _2980_/A vssd1 vssd1 vccd1 vccd1 _3129_/A sky130_fd_sc_hd__clkbuf_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _5314_/Q _4649_/X _4662_/S vssd1 vssd1 vccd1 vccd1 _4651_/B sky130_fd_sc_hd__mux2_1
X_3601_ _3780_/S vssd1 vssd1 vccd1 vccd1 _3767_/A sky130_fd_sc_hd__clkbuf_2
Xinput21 la1_data_in[11] vssd1 vssd1 vccd1 vccd1 _5338_/D sky130_fd_sc_hd__clkbuf_1
Xinput10 io_in[22] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_1
Xinput32 la1_data_in[21] vssd1 vssd1 vccd1 vccd1 _5348_/D sky130_fd_sc_hd__clkbuf_1
Xinput43 la1_data_in[6] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_2
X_4581_ _5300_/Q _4581_/B vssd1 vssd1 vccd1 vccd1 _4581_/X sky130_fd_sc_hd__or2_1
X_3532_ _3532_/A _3667_/A vssd1 vssd1 vccd1 vccd1 _3533_/B sky130_fd_sc_hd__nand2_1
X_3463_ _3464_/A _3464_/B vssd1 vssd1 vccd1 vccd1 _3465_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5202_ _5369_/CLK _5202_/D vssd1 vssd1 vccd1 vccd1 _5202_/Q sky130_fd_sc_hd__dfxtp_1
X_3394_ _3267_/X _3392_/Y _3393_/Y _3370_/X vssd1 vssd1 vccd1 vccd1 _3394_/X sky130_fd_sc_hd__a211o_1
X_5133_ _5313_/CLK _5133_/D vssd1 vssd1 vccd1 vccd1 _5133_/Q sky130_fd_sc_hd__dfxtp_1
X_5064_ _5064_/CLK _5064_/D vssd1 vssd1 vccd1 vccd1 _5064_/Q sky130_fd_sc_hd__dfxtp_1
X_4015_ _5124_/Q input11/X _4019_/S vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4917_ _4917_/A vssd1 vssd1 vccd1 vccd1 _5424_/D sky130_fd_sc_hd__clkbuf_1
X_4848_ _5373_/D _4840_/X _4847_/Y _4842_/X vssd1 vssd1 vccd1 vccd1 _5405_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4779_ _4783_/C _4779_/B vssd1 vssd1 vccd1 vccd1 _5366_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2963_ _2960_/X _2961_/Y _2962_/Y _3090_/A vssd1 vssd1 vccd1 vccd1 _2964_/B sky130_fd_sc_hd__a2bb2o_1
X_4702_ _4693_/A _4693_/B _4698_/X _5328_/Q vssd1 vssd1 vccd1 vccd1 _4702_/X sky130_fd_sc_hd__a31o_1
XFILLER_8_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2894_ _5376_/Q _5379_/Q _5378_/Q vssd1 vssd1 vccd1 vccd1 _2906_/A sky130_fd_sc_hd__or3_2
XFILLER_30_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633_ _4633_/A vssd1 vssd1 vccd1 vccd1 _5310_/D sky130_fd_sc_hd__clkbuf_1
X_4564_ _5293_/Q _4564_/B vssd1 vssd1 vccd1 vccd1 _4564_/X sky130_fd_sc_hd__or2_1
X_3515_ _5248_/Q _3673_/B vssd1 vssd1 vccd1 vccd1 _3532_/A sky130_fd_sc_hd__nor2_1
X_4495_ _5267_/Q _5105_/Q _4519_/S vssd1 vssd1 vccd1 vccd1 _4496_/A sky130_fd_sc_hd__mux2_1
X_3446_ _3853_/A _3841_/B _3446_/C _3446_/D vssd1 vssd1 vccd1 vccd1 _3447_/A sky130_fd_sc_hd__or4_1
X_3377_ _3377_/A _3419_/B vssd1 vssd1 vccd1 vccd1 _3378_/B sky130_fd_sc_hd__nand2_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5116_ _5116_/CLK _5116_/D vssd1 vssd1 vccd1 vccd1 _5116_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5047_ _5051_/CLK _5047_/D vssd1 vssd1 vccd1 vccd1 _5047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3300_ _3300_/A _3300_/B vssd1 vssd1 vccd1 vccd1 _3314_/A sky130_fd_sc_hd__xnor2_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4280_ _4280_/A vssd1 vssd1 vccd1 vccd1 _5211_/D sky130_fd_sc_hd__clkbuf_1
X_3231_ _5439_/Q _3197_/A _3229_/B _3229_/C _3230_/Y vssd1 vssd1 vccd1 vccd1 _3231_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _3163_/A _3163_/B vssd1 vssd1 vccd1 vccd1 _3181_/A sky130_fd_sc_hd__or2_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3093_ _3647_/A _5396_/Q _3139_/A vssd1 vssd1 vccd1 vccd1 _3097_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2946_ _2991_/A _5229_/Q vssd1 vssd1 vccd1 vccd1 _2946_/X sky130_fd_sc_hd__or2_1
X_2877_ _2867_/X _2871_/X _2876_/X _2854_/Y vssd1 vssd1 vccd1 vccd1 _2878_/B sky130_fd_sc_hd__o22a_1
X_4616_ _5289_/Q _5259_/Q _4616_/S vssd1 vssd1 vccd1 vccd1 _4616_/X sky130_fd_sc_hd__mux2_1
X_5596_ _5596_/A _2627_/Y vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__ebufn_8
X_4547_ _5287_/Q _5434_/Q _4549_/S vssd1 vssd1 vccd1 vccd1 _4548_/A sky130_fd_sc_hd__mux2_1
X_4478_ _4478_/A vssd1 vssd1 vccd1 vccd1 _5259_/D sky130_fd_sc_hd__clkbuf_1
X_3429_ _3396_/Y _3408_/A _3553_/A _3419_/B vssd1 vssd1 vccd1 vccd1 _3429_/X sky130_fd_sc_hd__a22o_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5484__74 vssd1 vssd1 vccd1 vccd1 _5484__74/HI _5562_/A sky130_fd_sc_hd__conb_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3780_ _3779_/X _5032_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3781_/A sky130_fd_sc_hd__mux2_1
X_2800_ _5127_/Q vssd1 vssd1 vccd1 vccd1 _2875_/S sky130_fd_sc_hd__clkbuf_2
X_2731_ _3764_/S vssd1 vssd1 vccd1 vccd1 _3726_/A sky130_fd_sc_hd__buf_2
XFILLER_13_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5450_ _5403_/Q _5450_/D vssd1 vssd1 vccd1 vccd1 _5603_/A sky130_fd_sc_hd__dfxtp_4
X_2662_ _2665_/A vssd1 vssd1 vccd1 vccd1 _2662_/Y sky130_fd_sc_hd__inv_2
X_4401_ _5237_/Q _4383_/X _4400_/X _4397_/X vssd1 vssd1 vccd1 vccd1 _5237_/D sky130_fd_sc_hd__o211a_1
X_2593_ _2597_/A vssd1 vssd1 vccd1 vccd1 _2593_/Y sky130_fd_sc_hd__inv_2
X_5381_ _5403_/Q _5381_/D vssd1 vssd1 vccd1 vccd1 _5381_/Q sky130_fd_sc_hd__dfxtp_4
X_4332_ _5325_/Q _5324_/Q vssd1 vssd1 vccd1 vccd1 _4586_/D sky130_fd_sc_hd__nor2_1
X_4263_ _4449_/C _4434_/B _3658_/B _3534_/B vssd1 vssd1 vccd1 vccd1 _4275_/A sky130_fd_sc_hd__a31o_1
X_3214_ _4992_/Q vssd1 vssd1 vccd1 vccd1 _3260_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4194_ _4193_/X _5187_/Q _4197_/S vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__mux2_1
X_3145_ _3081_/A _3081_/B _3081_/C _3102_/C _3144_/X vssd1 vssd1 vccd1 vccd1 _3150_/A
+ sky130_fd_sc_hd__a2111o_1
XFILLER_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3076_ _3076_/A vssd1 vssd1 vccd1 vccd1 _3076_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ _5099_/Q _3976_/X _3973_/X _4833_/A vssd1 vssd1 vccd1 vccd1 _5099_/D sky130_fd_sc_hd__a22o_1
X_2929_ _5372_/Q _2929_/B _2977_/C vssd1 vssd1 vccd1 vccd1 _2929_/X sky130_fd_sc_hd__or3_1
XFILLER_136_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5579_ _5579_/A _2606_/Y vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__ebufn_8
XFILLER_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput8 io_in[18] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4950_ _4953_/B _4953_/C _4094_/X vssd1 vssd1 vccd1 vccd1 _4950_/Y sky130_fd_sc_hd__a21oi_1
X_4881_ _4888_/C _4880_/Y _4841_/B vssd1 vssd1 vccd1 vccd1 _4881_/Y sky130_fd_sc_hd__o21ai_1
X_3901_ _5078_/Q _3898_/X _3956_/S vssd1 vssd1 vccd1 vccd1 _3902_/A sky130_fd_sc_hd__mux2_1
XFILLER_60_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3832_ _3835_/B _3835_/C vssd1 vssd1 vccd1 vccd1 _3834_/A sky130_fd_sc_hd__and2_1
XFILLER_20_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3763_ _3763_/A vssd1 vssd1 vccd1 vccd1 _5027_/D sky130_fd_sc_hd__clkbuf_1
X_2714_ _2714_/A vssd1 vssd1 vccd1 vccd1 _5036_/D sky130_fd_sc_hd__clkbuf_1
X_3694_ _3899_/B vssd1 vssd1 vccd1 vccd1 _4347_/S sky130_fd_sc_hd__buf_2
XFILLER_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5433_ _5435_/CLK _5433_/D vssd1 vssd1 vccd1 vccd1 _5433_/Q sky130_fd_sc_hd__dfxtp_1
X_2645_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2645_/Y sky130_fd_sc_hd__inv_2
X_5364_ _5371_/CLK _5364_/D vssd1 vssd1 vccd1 vccd1 _5364_/Q sky130_fd_sc_hd__dfxtp_1
X_2576_ _2578_/A vssd1 vssd1 vccd1 vccd1 _2576_/Y sky130_fd_sc_hd__inv_2
X_4315_ _4315_/A vssd1 vssd1 vccd1 vccd1 _5219_/D sky130_fd_sc_hd__clkbuf_1
X_5295_ _5437_/CLK _5295_/D vssd1 vssd1 vccd1 vccd1 _5295_/Q sky130_fd_sc_hd__dfxtp_1
X_4246_ _4252_/A _4246_/B vssd1 vssd1 vccd1 vccd1 _4247_/A sky130_fd_sc_hd__and2_1
X_4177_ _4176_/X _5182_/Q _4180_/S vssd1 vssd1 vccd1 vccd1 _4178_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3128_ _3074_/A _5383_/Q _3076_/A _5314_/Q vssd1 vssd1 vccd1 vccd1 _3129_/B sky130_fd_sc_hd__a22o_1
XFILLER_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3059_ _3134_/A _3059_/B vssd1 vssd1 vccd1 vccd1 _3060_/B sky130_fd_sc_hd__xor2_2
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_136_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5455__124 vssd1 vssd1 vccd1 vccd1 _5630_/A _5455__124/LO sky130_fd_sc_hd__conb_1
XFILLER_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4100_ _4100_/A _4100_/B vssd1 vssd1 vccd1 vccd1 _5156_/D sky130_fd_sc_hd__nor2_1
X_5080_ _5431_/CLK _5080_/D vssd1 vssd1 vccd1 vccd1 _5080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4031_ _2753_/A _3464_/B _4030_/Y vssd1 vssd1 vccd1 vccd1 _4041_/B sky130_fd_sc_hd__a21oi_1
XFILLER_52_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4933_ _4933_/A vssd1 vssd1 vccd1 vccd1 _5431_/D sky130_fd_sc_hd__clkbuf_1
X_4864_ _5408_/Q _5409_/Q _4864_/C vssd1 vssd1 vccd1 vccd1 _4869_/B sky130_fd_sc_hd__and3_1
XANTENNA_13 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 _3746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3815_ _3818_/C _3815_/B vssd1 vssd1 vccd1 vccd1 _5049_/D sky130_fd_sc_hd__nor2_1
XANTENNA_35 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4795_ _2942_/X _5388_/Q _4801_/S vssd1 vssd1 vccd1 vccd1 _4796_/A sky130_fd_sc_hd__mux2_1
X_3746_ _3746_/A0 _3746_/A1 _3764_/S vssd1 vssd1 vccd1 vccd1 _3746_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5416_ _5403_/Q _5416_/D vssd1 vssd1 vccd1 vccd1 _5416_/Q sky130_fd_sc_hd__dfxtp_1
X_3677_ _4115_/A _3677_/B vssd1 vssd1 vccd1 vccd1 _4292_/A sky130_fd_sc_hd__or2_1
X_2628_ _2628_/A vssd1 vssd1 vccd1 vccd1 _2628_/Y sky130_fd_sc_hd__inv_2
X_5347_ _5351_/CLK _5347_/D vssd1 vssd1 vccd1 vccd1 _5347_/Q sky130_fd_sc_hd__dfxtp_1
X_2559_ _5110_/Q vssd1 vssd1 vccd1 vccd1 _3705_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5278_ _5430_/CLK _5278_/D vssd1 vssd1 vccd1 vccd1 _5278_/Q sky130_fd_sc_hd__dfxtp_1
X_4229_ _4235_/A _4229_/B vssd1 vssd1 vccd1 vccd1 _4230_/A sky130_fd_sc_hd__and2_1
XFILLER_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4580_ _5295_/Q _4566_/A _4579_/X _4571_/X vssd1 vssd1 vccd1 vccd1 _5299_/D sky130_fd_sc_hd__o211a_1
X_3600_ _4115_/A _3604_/B _3733_/B vssd1 vssd1 vccd1 vccd1 _3780_/S sky130_fd_sc_hd__or3b_4
Xinput11 io_in[23] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
Xinput22 la1_data_in[12] vssd1 vssd1 vccd1 vccd1 _5339_/D sky130_fd_sc_hd__clkbuf_1
Xinput33 la1_data_in[22] vssd1 vssd1 vccd1 vccd1 _5349_/D sky130_fd_sc_hd__clkbuf_1
Xinput44 la1_data_in[7] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_2
X_3531_ _3531_/A vssd1 vssd1 vccd1 vccd1 _3667_/A sky130_fd_sc_hd__buf_2
XFILLER_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3462_ _3464_/B _3462_/B vssd1 vssd1 vccd1 vccd1 _3472_/A sky130_fd_sc_hd__or2_1
X_3393_ _3393_/A _3393_/B vssd1 vssd1 vccd1 vccd1 _3393_/Y sky130_fd_sc_hd__nand2_1
X_5201_ _5445_/CLK _5201_/D vssd1 vssd1 vccd1 vccd1 _5201_/Q sky130_fd_sc_hd__dfxtp_1
X_5132_ _5132_/CLK _5132_/D vssd1 vssd1 vccd1 vccd1 _5132_/Q sky130_fd_sc_hd__dfxtp_1
X_5063_ _5443_/CLK _5063_/D vssd1 vssd1 vccd1 vccd1 _5063_/Q sky130_fd_sc_hd__dfxtp_1
X_4014_ _4014_/A vssd1 vssd1 vccd1 vccd1 _5123_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4916_ _5424_/Q _2903_/B _4916_/S vssd1 vssd1 vccd1 vccd1 _4917_/A sky130_fd_sc_hd__mux2_1
X_4847_ _4901_/A _4847_/B vssd1 vssd1 vccd1 vccd1 _4847_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4778_ _5366_/Q _4780_/C _4742_/X vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__o21ai_1
X_3729_ _3729_/A _3729_/B _3729_/C vssd1 vssd1 vccd1 vccd1 _3729_/X sky130_fd_sc_hd__and3_1
XFILLER_29_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5032_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2962_ _2962_/A _2962_/B vssd1 vssd1 vccd1 vccd1 _2962_/Y sky130_fd_sc_hd__nor2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _4701_/A vssd1 vssd1 vccd1 vccd1 _5327_/D sky130_fd_sc_hd__clkbuf_1
X_2893_ _5303_/Q _2974_/A _2975_/A vssd1 vssd1 vccd1 vccd1 _2893_/X sky130_fd_sc_hd__a21o_1
X_4632_ _4632_/A _4632_/B vssd1 vssd1 vccd1 vccd1 _4633_/A sky130_fd_sc_hd__and2_1
XFILLER_8_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4563_ input5/X _4552_/X _4562_/X _4558_/X vssd1 vssd1 vccd1 vccd1 _5292_/D sky130_fd_sc_hd__o211a_1
X_4494_ _4532_/A vssd1 vssd1 vccd1 vccd1 _4519_/S sky130_fd_sc_hd__buf_2
X_3514_ _5004_/Q _5005_/Q _5006_/Q vssd1 vssd1 vccd1 vccd1 _3531_/A sky130_fd_sc_hd__or3b_1
X_3445_ _3823_/A _3835_/B _3445_/C vssd1 vssd1 vccd1 vccd1 _3446_/D sky130_fd_sc_hd__or3_1
X_3376_ _3551_/B vssd1 vssd1 vccd1 vccd1 _3563_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5115_/CLK _5115_/D vssd1 vssd1 vccd1 vccd1 _5115_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5046_ _5051_/CLK _5046_/D vssd1 vssd1 vccd1 vccd1 _5046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3823_/D _3284_/A vssd1 vssd1 vccd1 vccd1 _3230_/Y sky130_fd_sc_hd__nand2_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _3652_/A _3161_/B vssd1 vssd1 vccd1 vccd1 _3163_/B sky130_fd_sc_hd__xnor2_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3092_ _3126_/A vssd1 vssd1 vccd1 vccd1 _3647_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3994_ _4000_/A vssd1 vssd1 vccd1 vccd1 _3994_/X sky130_fd_sc_hd__buf_1
X_2945_ _5243_/Q vssd1 vssd1 vccd1 vccd1 _2991_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_136_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2876_ _2872_/X _2873_/X _2874_/X _2875_/X _2870_/A _3464_/A vssd1 vssd1 vccd1 vccd1
+ _2876_/X sky130_fd_sc_hd__mux4_1
X_5595_ _5595_/A _2626_/Y vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__ebufn_8
X_4615_ _4615_/A vssd1 vssd1 vccd1 vccd1 _5306_/D sky130_fd_sc_hd__clkbuf_1
X_4546_ _4546_/A vssd1 vssd1 vccd1 vccd1 _5286_/D sky130_fd_sc_hd__clkbuf_1
X_4477_ _5259_/Q _5097_/Q _4481_/S vssd1 vssd1 vccd1 vccd1 _4478_/A sky130_fd_sc_hd__mux2_1
X_3428_ _3709_/B _3428_/B vssd1 vssd1 vccd1 vccd1 _4075_/B sky130_fd_sc_hd__nand2_2
X_3359_ _3350_/S _3357_/X _3418_/S _3344_/X vssd1 vssd1 vccd1 vccd1 _3359_/X sky130_fd_sc_hd__a211o_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5029_ _5058_/CLK _5029_/D vssd1 vssd1 vccd1 vccd1 _5029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2730_ _3752_/A vssd1 vssd1 vccd1 vccd1 _3764_/S sky130_fd_sc_hd__clkbuf_2
X_2661_ _2665_/A vssd1 vssd1 vccd1 vccd1 _2661_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4400_ _4400_/A _4400_/B vssd1 vssd1 vccd1 vccd1 _4400_/X sky130_fd_sc_hd__or2_1
X_2592_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2597_/A sky130_fd_sc_hd__buf_2
X_5380_ _5403_/Q _5380_/D vssd1 vssd1 vccd1 vccd1 _5380_/Q sky130_fd_sc_hd__dfxtp_4
X_4331_ _5326_/Q vssd1 vssd1 vccd1 vccd1 _4586_/C sky130_fd_sc_hd__inv_2
X_4262_ _4262_/A vssd1 vssd1 vccd1 vccd1 _5207_/D sky130_fd_sc_hd__clkbuf_1
X_3213_ _3328_/A _3260_/D vssd1 vssd1 vccd1 vccd1 _3213_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4193_ _5411_/Q _5362_/Q _4199_/S vssd1 vssd1 vccd1 vccd1 _4193_/X sky130_fd_sc_hd__mux2_1
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3144_ _3146_/B _3144_/B _3132_/X vssd1 vssd1 vccd1 vccd1 _3144_/X sky130_fd_sc_hd__or3b_1
XFILLER_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3075_ _5240_/Q _3075_/B vssd1 vssd1 vccd1 vccd1 _3076_/A sky130_fd_sc_hd__and2_2
XFILLER_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3977_ _5098_/Q _3976_/X _3973_/X _4832_/B vssd1 vssd1 vccd1 vccd1 _5098_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2928_ _5238_/Q _2928_/B vssd1 vssd1 vccd1 vccd1 _2948_/A sky130_fd_sc_hd__xnor2_1
XFILLER_40_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2859_ _5016_/Q _5015_/Q _2859_/S vssd1 vssd1 vccd1 vccd1 _2859_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5578_ _5578_/A _2605_/Y vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__ebufn_8
X_4529_ _4529_/A vssd1 vssd1 vccd1 vccd1 _5278_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput9 io_in[19] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4880_ _5413_/Q _4880_/B vssd1 vssd1 vccd1 vccd1 _4880_/Y sky130_fd_sc_hd__nor2_1
X_3900_ _3959_/S vssd1 vssd1 vccd1 vccd1 _3956_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_32_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3831_ _3835_/C _3831_/B vssd1 vssd1 vccd1 vccd1 _5053_/D sky130_fd_sc_hd__nor2_1
X_3762_ _3761_/X _5027_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3763_/A sky130_fd_sc_hd__mux2_1
XFILLER_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2713_ _4348_/A _2713_/B vssd1 vssd1 vccd1 vccd1 _2714_/A sky130_fd_sc_hd__or2_1
X_3693_ _4589_/A _3693_/B vssd1 vssd1 vccd1 vccd1 _3899_/B sky130_fd_sc_hd__nor2_1
X_5432_ _5435_/CLK _5432_/D vssd1 vssd1 vccd1 vccd1 _5432_/Q sky130_fd_sc_hd__dfxtp_1
X_2644_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2644_/Y sky130_fd_sc_hd__inv_2
X_5363_ _5371_/CLK _5363_/D vssd1 vssd1 vccd1 vccd1 _5363_/Q sky130_fd_sc_hd__dfxtp_1
X_2575_ _2578_/A vssd1 vssd1 vccd1 vccd1 _2575_/Y sky130_fd_sc_hd__inv_2
X_4314_ _4313_/X _5219_/Q _4324_/S vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__mux2_1
X_5294_ _5437_/CLK _5294_/D vssd1 vssd1 vccd1 vccd1 _5294_/Q sky130_fd_sc_hd__dfxtp_1
X_4245_ _5202_/Q _5198_/Q _4251_/S vssd1 vssd1 vccd1 vccd1 _4246_/B sky130_fd_sc_hd__mux2_1
X_4176_ _5406_/Q _5357_/Q _4182_/S vssd1 vssd1 vccd1 vccd1 _4176_/X sky130_fd_sc_hd__mux2_1
X_3127_ _3126_/A _5398_/Q _3139_/A vssd1 vssd1 vccd1 vccd1 _3132_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3058_ _2994_/A _3056_/X _3066_/C vssd1 vssd1 vccd1 vccd1 _3059_/B sky130_fd_sc_hd__a21bo_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4030_ _4827_/A _5120_/Q vssd1 vssd1 vccd1 vccd1 _4030_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4932_ _5431_/Q _5382_/Q _4938_/S vssd1 vssd1 vccd1 vccd1 _4933_/A sky130_fd_sc_hd__mux2_1
XFILLER_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4863_ _4884_/A vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_14 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_25 _3746_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3814_ _5049_/Q _3813_/B _3800_/X vssd1 vssd1 vccd1 vccd1 _3815_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_36 _5589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4794_ _4794_/A vssd1 vssd1 vccd1 vccd1 _5387_/D sky130_fd_sc_hd__clkbuf_1
X_3745_ _3406_/Y _3427_/A _3751_/B _3427_/B vssd1 vssd1 vccd1 vccd1 _3745_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_137_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5415_ _5403_/Q _5415_/D vssd1 vssd1 vccd1 vccd1 _5415_/Q sky130_fd_sc_hd__dfxtp_1
X_3676_ _3676_/A vssd1 vssd1 vccd1 vccd1 _5006_/D sky130_fd_sc_hd__clkbuf_1
X_2627_ _2628_/A vssd1 vssd1 vccd1 vccd1 _2627_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5353_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5346_ _5351_/CLK _5346_/D vssd1 vssd1 vccd1 vccd1 _5346_/Q sky130_fd_sc_hd__dfxtp_1
X_2558_ _2558_/A _2558_/B vssd1 vssd1 vccd1 vccd1 _5112_/D sky130_fd_sc_hd__nor2_1
X_5277_ _5430_/CLK _5277_/D vssd1 vssd1 vccd1 vccd1 _5277_/Q sky130_fd_sc_hd__dfxtp_1
X_4228_ _5197_/Q input8/X _4234_/S vssd1 vssd1 vccd1 vccd1 _4229_/B sky130_fd_sc_hd__mux2_1
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4159_ _3665_/A _4421_/S _4165_/B vssd1 vssd1 vccd1 vccd1 _4161_/B sky130_fd_sc_hd__a21o_1
XFILLER_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 io_in[24] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 la1_data_in[13] vssd1 vssd1 vccd1 vccd1 _5340_/D sky130_fd_sc_hd__clkbuf_1
Xinput34 la1_data_in[23] vssd1 vssd1 vccd1 vccd1 _5350_/D sky130_fd_sc_hd__clkbuf_1
Xinput45 la1_data_in[8] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_2
X_3530_ _5220_/Q _3547_/B vssd1 vssd1 vccd1 vccd1 _3530_/X sky130_fd_sc_hd__or2_1
XFILLER_6_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3461_ _3461_/A vssd1 vssd1 vccd1 vccd1 _3464_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3392_ _3352_/S _3391_/X _3340_/Y vssd1 vssd1 vccd1 vccd1 _3392_/Y sky130_fd_sc_hd__o21ai_1
X_5200_ _5369_/CLK _5200_/D vssd1 vssd1 vccd1 vccd1 _5200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5131_ _5132_/CLK _5131_/D vssd1 vssd1 vccd1 vccd1 _5131_/Q sky130_fd_sc_hd__dfxtp_1
X_5062_ _5443_/CLK _5062_/D vssd1 vssd1 vccd1 vccd1 _5062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4013_ _5123_/Q input10/X _4019_/S vssd1 vssd1 vccd1 vccd1 _4014_/A sky130_fd_sc_hd__mux2_1
XFILLER_38_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4915_ _4915_/A vssd1 vssd1 vccd1 vccd1 _5423_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ _5404_/Q _5405_/Q vssd1 vssd1 vccd1 vccd1 _4847_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4777_ _5366_/Q _4780_/C vssd1 vssd1 vccd1 vccd1 _4783_/C sky130_fd_sc_hd__and2_1
X_3728_ _3728_/A1 _3734_/B _3726_/B vssd1 vssd1 vccd1 vccd1 _3729_/C sky130_fd_sc_hd__a21o_1
X_3659_ _4708_/A _3659_/B vssd1 vssd1 vccd1 vccd1 _3675_/S sky130_fd_sc_hd__or2_1
X_5329_ _5335_/CLK _5329_/D vssd1 vssd1 vccd1 vccd1 _5329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2961_ _2961_/A _2961_/B vssd1 vssd1 vccd1 vccd1 _2961_/Y sky130_fd_sc_hd__nor2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _4789_/B _4700_/B _4700_/C vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__and3_1
XFILLER_8_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2892_ _2892_/A vssd1 vssd1 vccd1 vccd1 _2975_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4631_ _5310_/Q _4630_/X _4640_/S vssd1 vssd1 vccd1 vccd1 _4632_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4562_ _5292_/Q _4564_/B vssd1 vssd1 vccd1 vccd1 _4562_/X sky130_fd_sc_hd__or2_1
XFILLER_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3513_ _4730_/B vssd1 vssd1 vccd1 vccd1 _4220_/C sky130_fd_sc_hd__clkbuf_2
X_4493_ _4493_/A vssd1 vssd1 vccd1 vccd1 _5266_/D sky130_fd_sc_hd__clkbuf_1
X_3444_ _3851_/A _3847_/B vssd1 vssd1 vccd1 vccd1 _3446_/C sky130_fd_sc_hd__nand2_1
X_3375_ _3370_/X _3373_/X _3374_/X _3267_/X _3393_/A vssd1 vssd1 vccd1 vccd1 _3387_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5114_ _5114_/CLK _5114_/D vssd1 vssd1 vccd1 vccd1 _5114_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5051_/CLK _5045_/D vssd1 vssd1 vccd1 vccd1 _5045_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4829_ _5419_/D _4720_/C _4829_/S vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3176_/A _3160_/B vssd1 vssd1 vccd1 vccd1 _3161_/B sky130_fd_sc_hd__and2_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ _3126_/A _3126_/B _5396_/Q vssd1 vssd1 vccd1 vccd1 _3097_/A sky130_fd_sc_hd__and3_1
XFILLER_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3993_ _3993_/A vssd1 vssd1 vccd1 vccd1 _5109_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2944_ _3120_/A vssd1 vssd1 vccd1 vccd1 _2944_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2875_ _5024_/Q _5023_/Q _2875_/S vssd1 vssd1 vccd1 vccd1 _2875_/X sky130_fd_sc_hd__mux2_1
X_4614_ _4632_/A _4614_/B vssd1 vssd1 vccd1 vccd1 _4615_/A sky130_fd_sc_hd__and2_1
X_5594_ _5594_/A _2625_/Y vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__ebufn_8
X_4545_ _5286_/Q _5433_/Q _4549_/S vssd1 vssd1 vccd1 vccd1 _4546_/A sky130_fd_sc_hd__mux2_1
X_4476_ _4476_/A vssd1 vssd1 vccd1 vccd1 _5258_/D sky130_fd_sc_hd__clkbuf_1
X_3427_ _3427_/A _3427_/B vssd1 vssd1 vccd1 vccd1 _3428_/B sky130_fd_sc_hd__nand2_1
X_3358_ _3358_/A vssd1 vssd1 vccd1 vccd1 _3418_/S sky130_fd_sc_hd__buf_4
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3289_ _3300_/A _3300_/B _3290_/C vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__a21oi_1
X_5028_ _5058_/CLK _5028_/D vssd1 vssd1 vccd1 vccd1 _5028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5475__65 vssd1 vssd1 vccd1 vccd1 _5475__65/HI _5552_/A sky130_fd_sc_hd__conb_1
XFILLER_29_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2660_ _2666_/A vssd1 vssd1 vccd1 vccd1 _2665_/A sky130_fd_sc_hd__buf_12
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2591_ _2591_/A vssd1 vssd1 vccd1 vccd1 _2591_/Y sky130_fd_sc_hd__inv_2
X_4330_ _5326_/Q _4692_/B _4333_/B vssd1 vssd1 vccd1 vccd1 _4330_/X sky130_fd_sc_hd__or3_1
X_4261_ _4789_/A _5207_/Q _4261_/S vssd1 vssd1 vccd1 vccd1 _4262_/A sky130_fd_sc_hd__mux2_1
X_3212_ _3295_/B _3292_/A _4990_/Q _4991_/Q vssd1 vssd1 vccd1 vccd1 _3260_/D sky130_fd_sc_hd__o211ai_2
X_4192_ _4192_/A vssd1 vssd1 vccd1 vccd1 _5186_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3143_ _3148_/A _3148_/B vssd1 vssd1 vccd1 vccd1 _3166_/A sky130_fd_sc_hd__or2_1
XFILLER_39_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3074_ _3074_/A vssd1 vssd1 vccd1 vccd1 _3074_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3976_ _3983_/A vssd1 vssd1 vccd1 vccd1 _3976_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2927_ _2950_/A _5388_/Q vssd1 vssd1 vccd1 vccd1 _2928_/B sky130_fd_sc_hd__nand2_1
X_2858_ _5018_/Q _5017_/Q _2859_/S vssd1 vssd1 vccd1 vccd1 _2858_/X sky130_fd_sc_hd__mux2_1
X_5577_ _5577_/A _2603_/Y vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__ebufn_8
X_2789_ _5302_/Q _5150_/Q _2789_/C vssd1 vssd1 vccd1 vccd1 _3415_/A sky130_fd_sc_hd__and3_4
X_4528_ _5278_/Q _5425_/Q _4530_/S vssd1 vssd1 vccd1 vccd1 _4529_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4459_ _4450_/A _4445_/X _4455_/X _5253_/Q vssd1 vssd1 vccd1 vccd1 _4459_/X sky130_fd_sc_hd__a31o_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3830_ _3829_/A _3828_/A _3826_/X vssd1 vssd1 vccd1 vccd1 _3831_/B sky130_fd_sc_hd__o21ai_1
XFILLER_32_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3761_ _3750_/X _3759_/X _3760_/X _3754_/X vssd1 vssd1 vccd1 vccd1 _3761_/X sky130_fd_sc_hd__a22o_1
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2712_ _2706_/Y _3715_/A _3596_/A vssd1 vssd1 vccd1 vccd1 _2713_/B sky130_fd_sc_hd__o21a_1
XFILLER_9_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3692_ _4594_/A _3691_/Y _3625_/C _4594_/B vssd1 vssd1 vccd1 vccd1 _3693_/B sky130_fd_sc_hd__a211o_1
X_5431_ _5431_/CLK _5431_/D vssd1 vssd1 vccd1 vccd1 _5431_/Q sky130_fd_sc_hd__dfxtp_1
X_2643_ _2647_/A vssd1 vssd1 vccd1 vccd1 _2643_/Y sky130_fd_sc_hd__inv_2
X_5362_ _5371_/CLK _5362_/D vssd1 vssd1 vccd1 vccd1 _5362_/Q sky130_fd_sc_hd__dfxtp_1
X_2574_ _2578_/A vssd1 vssd1 vccd1 vccd1 _2574_/Y sky130_fd_sc_hd__inv_2
X_4313_ _5169_/Q _3537_/X _3674_/B _4311_/Y _4312_/X vssd1 vssd1 vccd1 vccd1 _4313_/X
+ sky130_fd_sc_hd__a221o_1
X_5293_ _5437_/CLK _5293_/D vssd1 vssd1 vccd1 vccd1 _5293_/Q sky130_fd_sc_hd__dfxtp_1
X_4244_ _4244_/A vssd1 vssd1 vccd1 vccd1 _5201_/D sky130_fd_sc_hd__clkbuf_1
X_4175_ _4175_/A vssd1 vssd1 vccd1 vccd1 _5181_/D sky130_fd_sc_hd__clkbuf_1
X_3999__7 _3999__7/A vssd1 vssd1 vccd1 vccd1 _5114_/CLK sky130_fd_sc_hd__inv_2
X_3126_ _3126_/A _3126_/B _5398_/Q vssd1 vssd1 vccd1 vccd1 _3132_/A sky130_fd_sc_hd__and3_1
XFILLER_28_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3057_ _3057_/A _3057_/B _3057_/C vssd1 vssd1 vccd1 vccd1 _3066_/C sky130_fd_sc_hd__or3_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ _5092_/Q _3958_/X _3959_/S vssd1 vssd1 vccd1 vccd1 _3960_/A sky130_fd_sc_hd__mux2_1
X_5629_ _5629_/A _2667_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__ebufn_8
XFILLER_19_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4931_ _4931_/A vssd1 vssd1 vccd1 vccd1 _5430_/D sky130_fd_sc_hd__clkbuf_1
X_4862_ _5376_/D _4840_/X _4859_/Y _4861_/X vssd1 vssd1 vccd1 vccd1 _5408_/D sky130_fd_sc_hd__o211a_1
XFILLER_60_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3813_ _5049_/Q _3813_/B vssd1 vssd1 vccd1 vccd1 _3818_/C sky130_fd_sc_hd__and2_1
XFILLER_20_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4793_ _2918_/X _5387_/Q _4801_/S vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__mux2_1
XANTENNA_26 _4348_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_15 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 _5590_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3744_ _3841_/A _3847_/A vssd1 vssd1 vccd1 vccd1 _3751_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3675_ _3674_/Y _5006_/Q _3675_/S vssd1 vssd1 vccd1 vccd1 _3676_/A sky130_fd_sc_hd__mux2_1
X_2626_ _2628_/A vssd1 vssd1 vccd1 vccd1 _2626_/Y sky130_fd_sc_hd__inv_2
X_5414_ _5403_/Q _5414_/D vssd1 vssd1 vccd1 vccd1 _5414_/Q sky130_fd_sc_hd__dfxtp_1
X_5345_ _5351_/CLK _5345_/D vssd1 vssd1 vccd1 vccd1 _5345_/Q sky130_fd_sc_hd__dfxtp_1
X_2557_ _2743_/A _2562_/A _2544_/X vssd1 vssd1 vccd1 vccd1 _2558_/B sky130_fd_sc_hd__o21ai_1
X_5276_ _5430_/CLK _5276_/D vssd1 vssd1 vccd1 vccd1 _5276_/Q sky130_fd_sc_hd__dfxtp_1
X_4227_ _4227_/A vssd1 vssd1 vccd1 vccd1 _5196_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4158_ _4158_/A _4433_/A vssd1 vssd1 vccd1 vccd1 _4165_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4089_ _5153_/Q _4086_/A _4088_/Y vssd1 vssd1 vccd1 vccd1 _5153_/D sky130_fd_sc_hd__o21a_1
X_3109_ _3126_/B _3109_/B vssd1 vssd1 vccd1 vccd1 _3114_/A sky130_fd_sc_hd__xnor2_1
XFILLER_24_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5526__116 vssd1 vssd1 vccd1 vccd1 _5526__116/HI _5526__116/LO sky130_fd_sc_hd__conb_1
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput13 io_in[25] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__clkbuf_1
Xinput24 la1_data_in[14] vssd1 vssd1 vccd1 vccd1 _5341_/D sky130_fd_sc_hd__clkbuf_1
Xinput35 la1_data_in[24] vssd1 vssd1 vccd1 vccd1 _5351_/D sky130_fd_sc_hd__clkbuf_1
Xinput46 la1_data_in[9] vssd1 vssd1 vccd1 vccd1 _4945_/C sky130_fd_sc_hd__buf_2
XFILLER_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3460_ _3448_/Y _3449_/Y _3451_/Y _3455_/X _3459_/Y vssd1 vssd1 vccd1 vccd1 _5589_/A
+ sky130_fd_sc_hd__a311oi_4
X_3391_ _3343_/A _3390_/Y _3372_/B vssd1 vssd1 vccd1 vccd1 _3391_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5130_ _5132_/CLK _5130_/D vssd1 vssd1 vccd1 vccd1 _5130_/Q sky130_fd_sc_hd__dfxtp_1
X_5061_ _5439_/CLK _5061_/D vssd1 vssd1 vccd1 vccd1 _5061_/Q sky130_fd_sc_hd__dfxtp_1
X_4012_ _4012_/A _5134_/D vssd1 vssd1 vccd1 vccd1 _4019_/S sky130_fd_sc_hd__nor2_8
X_4914_ _5423_/Q _2903_/C _4916_/S vssd1 vssd1 vccd1 vccd1 _4915_/A sky130_fd_sc_hd__mux2_1
X_4845_ _4884_/A vssd1 vssd1 vccd1 vccd1 _4901_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4776_ _4780_/C _4776_/B vssd1 vssd1 vccd1 vccd1 _5365_/D sky130_fd_sc_hd__nor2_1
X_3727_ _3710_/X _3726_/X _5020_/Q _4043_/A vssd1 vssd1 vccd1 vccd1 _5020_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_20_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3658_ _3658_/A _3658_/B vssd1 vssd1 vccd1 vccd1 _3659_/B sky130_fd_sc_hd__or2_1
X_2609_ _2609_/A vssd1 vssd1 vccd1 vccd1 _2609_/Y sky130_fd_sc_hd__inv_2
X_3589_ _5219_/Q _3529_/A _4434_/C _4355_/A vssd1 vssd1 vccd1 vccd1 _3589_/X sky130_fd_sc_hd__o211a_1
X_5328_ _5328_/CLK _5328_/D vssd1 vssd1 vccd1 vccd1 _5328_/Q sky130_fd_sc_hd__dfxtp_1
X_5259_ _5435_/CLK _5259_/D vssd1 vssd1 vccd1 vccd1 _5259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2960_ _2961_/A _2961_/B _3090_/A vssd1 vssd1 vccd1 vccd1 _2960_/X sky130_fd_sc_hd__a21o_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2891_ _5240_/Q vssd1 vssd1 vccd1 vccd1 _2892_/A sky130_fd_sc_hd__inv_2
XFILLER_8_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4630_ _5292_/Q _5262_/Q _4639_/S vssd1 vssd1 vccd1 vccd1 _4630_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4561_ input4/X _4552_/X _4560_/X _4558_/X vssd1 vssd1 vccd1 vccd1 _5291_/D sky130_fd_sc_hd__o211a_1
XFILLER_7_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3512_ _5247_/Q _5246_/Q vssd1 vssd1 vccd1 vccd1 _4730_/B sky130_fd_sc_hd__nor2_1
X_4492_ _5266_/Q _5104_/Q _4492_/S vssd1 vssd1 vccd1 vccd1 _4493_/A sky130_fd_sc_hd__mux2_1
X_3443_ _3824_/B _3824_/C _3841_/A vssd1 vssd1 vccd1 vccd1 _3847_/B sky130_fd_sc_hd__and3_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _3374_/A _3374_/B vssd1 vssd1 vccd1 vccd1 _3374_/X sky130_fd_sc_hd__or2_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _5113_/CLK _5113_/D vssd1 vssd1 vccd1 vccd1 _5113_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5044_ _5245_/CLK _5044_/D vssd1 vssd1 vccd1 vccd1 _5044_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4828_ _4828_/A vssd1 vssd1 vccd1 vccd1 _5419_/D sky130_fd_sc_hd__clkbuf_1
X_4759_ _5360_/Q _4757_/A _4746_/X vssd1 vssd1 vccd1 vccd1 _4760_/B sky130_fd_sc_hd__o21ai_1
XFILLER_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_12_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5328_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_17_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3090_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3646_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _4789_/A _4571_/A vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__and2_1
XFILLER_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2943_ _4791_/A _5233_/Q vssd1 vssd1 vccd1 vccd1 _3120_/A sky130_fd_sc_hd__nand2_1
X_2874_ _5026_/Q _5025_/Q _2875_/S vssd1 vssd1 vccd1 vccd1 _2874_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4613_ _5306_/Q _4612_/X _4617_/S vssd1 vssd1 vccd1 vccd1 _4614_/B sky130_fd_sc_hd__mux2_1
X_5593_ _5593_/A _2624_/Y vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__ebufn_8
X_4544_ _4544_/A vssd1 vssd1 vccd1 vccd1 _5285_/D sky130_fd_sc_hd__clkbuf_1
X_4475_ _5258_/Q _5096_/Q _4481_/S vssd1 vssd1 vccd1 vccd1 _4476_/A sky130_fd_sc_hd__mux2_1
X_3426_ _3427_/A _3427_/B vssd1 vssd1 vccd1 vccd1 _3709_/B sky130_fd_sc_hd__or2_1
X_3357_ _3357_/A vssd1 vssd1 vccd1 vccd1 _3357_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ _3409_/A _3287_/Y _3252_/S _3280_/Y vssd1 vssd1 vccd1 vccd1 _3290_/C sky130_fd_sc_hd__a2bb2o_1
X_5027_ _5032_/CLK _5027_/D vssd1 vssd1 vccd1 vccd1 _5027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2590_ _2591_/A vssd1 vssd1 vccd1 vccd1 _2590_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ _4260_/A vssd1 vssd1 vccd1 vccd1 _5206_/D sky130_fd_sc_hd__clkbuf_1
X_3211_ _3211_/A vssd1 vssd1 vccd1 vccd1 _3295_/B sky130_fd_sc_hd__clkbuf_2
X_4191_ _4190_/X _5186_/Q _4197_/S vssd1 vssd1 vccd1 vccd1 _4192_/A sky130_fd_sc_hd__mux2_1
X_3142_ _3142_/A _3142_/B vssd1 vssd1 vccd1 vccd1 _3148_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3073_ _3129_/A vssd1 vssd1 vccd1 vccd1 _3176_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3975_ _5097_/Q _3966_/X _3973_/X _4832_/A vssd1 vssd1 vccd1 vccd1 _5097_/D sky130_fd_sc_hd__a22o_1
X_2926_ _5234_/Q vssd1 vssd1 vccd1 vccd1 _3023_/A sky130_fd_sc_hd__buf_2
X_2857_ _2855_/X _2856_/X _2860_/S vssd1 vssd1 vccd1 vccd1 _2857_/X sky130_fd_sc_hd__mux2_1
XFILLER_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5576_ _5576_/A _2602_/Y vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__ebufn_8
X_2788_ _2788_/A vssd1 vssd1 vccd1 vccd1 _2789_/C sky130_fd_sc_hd__inv_2
X_4527_ _4527_/A vssd1 vssd1 vccd1 vccd1 _5277_/D sky130_fd_sc_hd__clkbuf_1
X_4458_ _4458_/A vssd1 vssd1 vccd1 vccd1 _5252_/D sky130_fd_sc_hd__clkbuf_1
X_3409_ _3409_/A _3553_/A _3409_/C vssd1 vssd1 vccd1 vccd1 _3409_/X sky130_fd_sc_hd__and3_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4389_ _5197_/Q _5167_/Q _4399_/S vssd1 vssd1 vccd1 vccd1 _4390_/B sky130_fd_sc_hd__mux2_1
XFILLER_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3760_ _3760_/A0 _3760_/A1 _3773_/S vssd1 vssd1 vccd1 vccd1 _3760_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2711_ _5036_/Q vssd1 vssd1 vccd1 vccd1 _3596_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5430_ _5430_/CLK _5430_/D vssd1 vssd1 vccd1 vccd1 _5430_/Q sky130_fd_sc_hd__dfxtp_1
X_3691_ _4328_/B _3945_/B vssd1 vssd1 vccd1 vccd1 _3691_/Y sky130_fd_sc_hd__nor2_1
X_2642_ _2666_/A vssd1 vssd1 vccd1 vccd1 _2647_/A sky130_fd_sc_hd__buf_2
X_5361_ _5444_/CLK _5361_/D vssd1 vssd1 vccd1 vccd1 _5361_/Q sky130_fd_sc_hd__dfxtp_1
X_2573_ _2698_/A vssd1 vssd1 vccd1 vccd1 _2578_/A sky130_fd_sc_hd__clkbuf_2
X_4312_ _5215_/Q _3543_/B _3535_/A vssd1 vssd1 vccd1 vccd1 _4312_/X sky130_fd_sc_hd__o21a_1
X_5292_ _5437_/CLK _5292_/D vssd1 vssd1 vccd1 vccd1 _5292_/Q sky130_fd_sc_hd__dfxtp_1
X_4243_ _4252_/A _4243_/B vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__and2_1
X_4174_ _4173_/X _5181_/Q _4180_/S vssd1 vssd1 vccd1 vccd1 _4175_/A sky130_fd_sc_hd__mux2_1
X_3125_ _3144_/B _3117_/B _3084_/A _3146_/A vssd1 vssd1 vccd1 vccd1 _3135_/A sky130_fd_sc_hd__o211a_1
XFILLER_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3056_ _3057_/A _3057_/B _3057_/C vssd1 vssd1 vccd1 vccd1 _3056_/X sky130_fd_sc_hd__o21a_1
XFILLER_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3958_ _5266_/Q _3915_/A _3943_/X _5088_/Q _3947_/X vssd1 vssd1 vccd1 vccd1 _3958_/X
+ sky130_fd_sc_hd__a221o_1
X_3889_ _3889_/A vssd1 vssd1 vccd1 vccd1 _5077_/D sky130_fd_sc_hd__clkbuf_1
X_2909_ _5237_/Q vssd1 vssd1 vccd1 vccd1 _2910_/A sky130_fd_sc_hd__inv_2
X_5628_ _5629_/A _2665_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__ebufn_8
X_5559_ _5559_/A _2583_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4930_ _5430_/Q _5381_/Q _4938_/S vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__mux2_1
X_4861_ _4861_/A vssd1 vssd1 vccd1 vccd1 _4861_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3812_ _3813_/B _3812_/B vssd1 vssd1 vccd1 vccd1 _5048_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_16 _5377_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4792_ _4825_/S vssd1 vssd1 vccd1 vccd1 _4801_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_27 _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3743_ _5024_/Q _3602_/X _3740_/X _3742_/X vssd1 vssd1 vccd1 vccd1 _5024_/D sky130_fd_sc_hd__a22o_1
X_3674_ _5006_/Q _3674_/B vssd1 vssd1 vccd1 vccd1 _3674_/Y sky130_fd_sc_hd__nor2_1
X_5413_ _5403_/Q _5413_/D vssd1 vssd1 vccd1 vccd1 _5413_/Q sky130_fd_sc_hd__dfxtp_1
X_2625_ _2628_/A vssd1 vssd1 vccd1 vccd1 _2625_/Y sky130_fd_sc_hd__inv_2
X_5344_ _5351_/CLK _5344_/D vssd1 vssd1 vccd1 vccd1 _5344_/Q sky130_fd_sc_hd__dfxtp_1
X_2556_ _2556_/A _2556_/B vssd1 vssd1 vccd1 vccd1 _5113_/D sky130_fd_sc_hd__nor2_1
X_5275_ _5430_/CLK _5275_/D vssd1 vssd1 vccd1 vccd1 _5275_/Q sky130_fd_sc_hd__dfxtp_1
X_4226_ _4235_/A _4226_/B vssd1 vssd1 vccd1 vccd1 _4227_/A sky130_fd_sc_hd__and2_1
X_4157_ _4154_/A _4155_/X _5354_/Q _4156_/Y vssd1 vssd1 vccd1 vccd1 _4433_/A sky130_fd_sc_hd__o211a_1
X_3108_ _3108_/A _5397_/Q vssd1 vssd1 vccd1 vccd1 _3109_/B sky130_fd_sc_hd__and2_1
X_4088_ _2781_/B _4092_/B _4954_/A vssd1 vssd1 vccd1 vccd1 _4088_/Y sky130_fd_sc_hd__a21oi_1
X_3039_ _3013_/C _3067_/B _3038_/X vssd1 vssd1 vccd1 vccd1 _3040_/B sky130_fd_sc_hd__o21a_1
XFILLER_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5505__95 vssd1 vssd1 vccd1 vccd1 _5505__95/HI _5608_/A sky130_fd_sc_hd__conb_1
XFILLER_47_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput14 io_in[26] vssd1 vssd1 vccd1 vccd1 _2786_/C sky130_fd_sc_hd__buf_2
Xinput25 la1_data_in[15] vssd1 vssd1 vccd1 vccd1 _5342_/D sky130_fd_sc_hd__clkbuf_1
Xinput36 la1_data_in[25] vssd1 vssd1 vccd1 vccd1 _5352_/D sky130_fd_sc_hd__clkbuf_1
X_3390_ _3390_/A _3390_/B vssd1 vssd1 vccd1 vccd1 _3390_/Y sky130_fd_sc_hd__nand2_1
X_5060_ _5439_/CLK _5060_/D vssd1 vssd1 vccd1 vccd1 _5060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4011_ _3705_/A _2752_/B _4010_/X _3750_/A vssd1 vssd1 vccd1 vccd1 _5134_/D sky130_fd_sc_hd__o31ai_4
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4913_ _4913_/A vssd1 vssd1 vccd1 vccd1 _5422_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4844_ _4844_/A vssd1 vssd1 vccd1 vccd1 _4884_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4775_ _5365_/Q _4773_/A _4762_/X vssd1 vssd1 vccd1 vccd1 _4776_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3726_ _3726_/A _3726_/B _3726_/C_N vssd1 vssd1 vccd1 vccd1 _3726_/X sky130_fd_sc_hd__or3b_1
X_3657_ _3645_/Y _2925_/X _3656_/Y _2944_/X vssd1 vssd1 vccd1 vccd1 _5003_/D sky130_fd_sc_hd__o22ai_1
X_2608_ _2609_/A vssd1 vssd1 vccd1 vccd1 _2608_/Y sky130_fd_sc_hd__inv_2
X_3588_ _4434_/A vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__clkbuf_2
X_5327_ _5328_/CLK _5327_/D vssd1 vssd1 vccd1 vccd1 _5327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2539_ _5114_/Q _2736_/B _2558_/A vssd1 vssd1 vccd1 vccd1 _2554_/A sky130_fd_sc_hd__and3_1
X_5258_ _5305_/CLK _5258_/D vssd1 vssd1 vccd1 vccd1 _5258_/Q sky130_fd_sc_hd__dfxtp_1
X_5189_ _5369_/CLK _5189_/D vssd1 vssd1 vccd1 vccd1 _5189_/Q sky130_fd_sc_hd__dfxtp_1
X_4209_ _4209_/A vssd1 vssd1 vccd1 vccd1 _5191_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_44_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_137_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2890_ _2890_/A vssd1 vssd1 vccd1 vccd1 _2974_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4560_ _5291_/Q _4564_/B vssd1 vssd1 vccd1 vccd1 _4560_/X sky130_fd_sc_hd__or2_1
XFILLER_8_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3511_ _3662_/C _3526_/A vssd1 vssd1 vccd1 vccd1 _3511_/Y sky130_fd_sc_hd__nor2_1
X_4491_ _4491_/A vssd1 vssd1 vccd1 vccd1 _5265_/D sky130_fd_sc_hd__clkbuf_1
X_3442_ _3442_/A vssd1 vssd1 vccd1 vccd1 _3841_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3373_ _3374_/A _3373_/B _3373_/C vssd1 vssd1 vccd1 vccd1 _3373_/X sky130_fd_sc_hd__or3_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5112_/CLK _5112_/D vssd1 vssd1 vccd1 vccd1 _5112_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5051_/CLK _5043_/D vssd1 vssd1 vccd1 vccd1 _5043_/Q sky130_fd_sc_hd__dfxtp_1
X_5496__86 vssd1 vssd1 vccd1 vccd1 _5496__86/HI _5592_/A sky130_fd_sc_hd__conb_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4827_ _4827_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _4828_/A sky130_fd_sc_hd__and2_1
XFILLER_21_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4758_ _5360_/Q _5359_/Q _4758_/C vssd1 vssd1 vccd1 vccd1 _4765_/C sky130_fd_sc_hd__and3_1
X_4689_ _4589_/Y _3946_/B _4586_/D _4694_/B vssd1 vssd1 vccd1 vccd1 _4689_/X sky130_fd_sc_hd__a211o_1
X_3709_ _3709_/A _3709_/B _5040_/Q vssd1 vssd1 vccd1 vccd1 _3736_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_3991_ _4203_/A vssd1 vssd1 vccd1 vccd1 _4789_/A sky130_fd_sc_hd__clkbuf_4
X_2942_ _4831_/B vssd1 vssd1 vccd1 vccd1 _2942_/X sky130_fd_sc_hd__clkbuf_4
X_2873_ _5028_/Q _5027_/Q _2875_/S vssd1 vssd1 vccd1 vccd1 _2873_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5592_ _5592_/A _2622_/Y vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__ebufn_8
X_4612_ input5/X _5258_/Q _4616_/S vssd1 vssd1 vccd1 vccd1 _4612_/X sky130_fd_sc_hd__mux2_1
X_4543_ _5285_/Q _5432_/Q _4549_/S vssd1 vssd1 vccd1 vccd1 _4544_/A sky130_fd_sc_hd__mux2_1
X_4474_ _4474_/A vssd1 vssd1 vccd1 vccd1 _5257_/D sky130_fd_sc_hd__clkbuf_1
X_3425_ _3853_/A _3824_/B _3749_/B vssd1 vssd1 vccd1 vccd1 _3427_/B sky130_fd_sc_hd__or3_1
X_3356_ _3356_/A _3356_/B vssd1 vssd1 vccd1 vccd1 _3393_/B sky130_fd_sc_hd__xnor2_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3287_ _3442_/A _3772_/B _3286_/C vssd1 vssd1 vccd1 vccd1 _3287_/Y sky130_fd_sc_hd__a21oi_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5032_/CLK _5026_/D vssd1 vssd1 vccd1 vccd1 _5026_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3210_ _3211_/A _3292_/A vssd1 vssd1 vccd1 vccd1 _3328_/A sky130_fd_sc_hd__or2_2
X_4190_ _5410_/Q _5361_/Q _4199_/S vssd1 vssd1 vccd1 vccd1 _4190_/X sky130_fd_sc_hd__mux2_1
X_3141_ _3176_/A _3141_/B vssd1 vssd1 vccd1 vccd1 _3142_/B sky130_fd_sc_hd__and2_1
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5466__56 vssd1 vssd1 vccd1 vccd1 _5466__56/HI _5543_/A sky130_fd_sc_hd__conb_1
XFILLER_54_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3072_ _3130_/A vssd1 vssd1 vccd1 vccd1 _3142_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3974_ _5096_/Q _3966_/X _3973_/X _2990_/X vssd1 vssd1 vccd1 vccd1 _5096_/D sky130_fd_sc_hd__a22o_1
X_2925_ _3027_/A vssd1 vssd1 vccd1 vccd1 _2925_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2856_ _5020_/Q _5019_/Q _2859_/S vssd1 vssd1 vccd1 vccd1 _2856_/X sky130_fd_sc_hd__mux2_1
X_5575_ _5575_/A _2601_/Y vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__ebufn_8
X_2787_ _5446_/Q _2787_/B _5445_/Q _5227_/Q vssd1 vssd1 vccd1 vccd1 _2788_/A sky130_fd_sc_hd__or4b_1
X_4526_ _5277_/Q _5424_/Q _4530_/S vssd1 vssd1 vccd1 vccd1 _4527_/A sky130_fd_sc_hd__mux2_1
X_4457_ _4789_/B _4457_/B _4457_/C vssd1 vssd1 vccd1 vccd1 _4458_/A sky130_fd_sc_hd__and3_1
X_3408_ _3408_/A _3408_/B vssd1 vssd1 vccd1 vccd1 _3409_/C sky130_fd_sc_hd__nor2_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4388_ _5233_/Q _4383_/X _4387_/X _4378_/X vssd1 vssd1 vccd1 vccd1 _5233_/D sky130_fd_sc_hd__o211a_1
X_3339_ _3390_/A _3390_/B _3343_/A vssd1 vssd1 vccd1 vccd1 _3340_/B sky130_fd_sc_hd__mux2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ _5339_/CLK _5009_/D vssd1 vssd1 vccd1 vccd1 _5009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5480__70 vssd1 vssd1 vccd1 vccd1 _5480__70/HI _5557_/A sky130_fd_sc_hd__conb_1
XFILLER_26_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2710_ _5110_/Q _3705_/D _2729_/C vssd1 vssd1 vccd1 vccd1 _3715_/A sky130_fd_sc_hd__or3_1
X_3690_ _5326_/Q _4692_/B _4333_/B vssd1 vssd1 vccd1 vccd1 _3945_/B sky130_fd_sc_hd__nor3_2
X_2641_ input1/X vssd1 vssd1 vccd1 vccd1 _2666_/A sky130_fd_sc_hd__buf_8
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5360_ _5444_/CLK _5360_/D vssd1 vssd1 vccd1 vccd1 _5360_/Q sky130_fd_sc_hd__dfxtp_1
X_2572_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2572_/Y sky130_fd_sc_hd__inv_2
X_5291_ _5437_/CLK _5291_/D vssd1 vssd1 vccd1 vccd1 _5291_/Q sky130_fd_sc_hd__dfxtp_1
X_4311_ _5207_/Q vssd1 vssd1 vccd1 vccd1 _4311_/Y sky130_fd_sc_hd__inv_2
X_4242_ _5201_/Q _5197_/Q _4251_/S vssd1 vssd1 vccd1 vccd1 _4243_/B sky130_fd_sc_hd__mux2_1
X_4173_ _5405_/Q _5356_/Q _4182_/S vssd1 vssd1 vccd1 vccd1 _4173_/X sky130_fd_sc_hd__mux2_1
X_3124_ _5382_/Q _3028_/X _4834_/B _3120_/X _3123_/X vssd1 vssd1 vccd1 vccd1 _5382_/D
+ sky130_fd_sc_hd__o221a_1
X_3055_ _3130_/A _3055_/B vssd1 vssd1 vccd1 vccd1 _3057_/C sky130_fd_sc_hd__xnor2_2
XFILLER_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3957_ _3957_/A vssd1 vssd1 vccd1 vccd1 _5091_/D sky130_fd_sc_hd__clkbuf_1
X_2908_ _5451_/Q _4975_/B _2905_/X _2907_/X vssd1 vssd1 vccd1 vccd1 _2908_/X sky130_fd_sc_hd__o211a_1
XFILLER_137_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3888_ hold16/A _4837_/B _3888_/S vssd1 vssd1 vccd1 vccd1 _3889_/A sky130_fd_sc_hd__mux2_1
XFILLER_137_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5627_ _5629_/A _2664_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[23] sky130_fd_sc_hd__ebufn_8
X_2839_ _5017_/Q _3474_/B vssd1 vssd1 vccd1 vccd1 _2839_/X sky130_fd_sc_hd__and2_1
X_5558_ _5558_/A _2582_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[24] sky130_fd_sc_hd__ebufn_8
X_4509_ _5271_/Q _4514_/B _4553_/A vssd1 vssd1 vccd1 vccd1 _4509_/X sky130_fd_sc_hd__or3b_1
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_7_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5064_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_2_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4860_ _4902_/A vssd1 vssd1 vccd1 vccd1 _4861_/A sky130_fd_sc_hd__clkbuf_2
X_3811_ _5048_/Q _3809_/A _3800_/X vssd1 vssd1 vccd1 vccd1 _3812_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_17 _5379_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4791_ _4791_/A _5232_/Q vssd1 vssd1 vccd1 vccd1 _4825_/S sky130_fd_sc_hd__nand2_2
XANTENNA_28 _4685_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3742_ _3742_/A1 _3734_/B _4075_/B _3741_/X vssd1 vssd1 vccd1 vccd1 _3742_/X sky130_fd_sc_hd__a22o_1
X_3673_ _4112_/A _3673_/B _4432_/A vssd1 vssd1 vccd1 vccd1 _3674_/B sky130_fd_sc_hd__and3_2
X_5412_ _5403_/Q _5412_/D vssd1 vssd1 vccd1 vccd1 _5412_/Q sky130_fd_sc_hd__dfxtp_1
X_2624_ _2628_/A vssd1 vssd1 vccd1 vccd1 _2624_/Y sky130_fd_sc_hd__inv_2
X_5343_ _5351_/CLK _5343_/D vssd1 vssd1 vccd1 vccd1 _5343_/Q sky130_fd_sc_hd__dfxtp_1
X_2555_ _2736_/B _2558_/A _2544_/X vssd1 vssd1 vccd1 vccd1 _2556_/B sky130_fd_sc_hd__o21ai_1
X_5274_ _5430_/CLK _5274_/D vssd1 vssd1 vccd1 vccd1 _5274_/Q sky130_fd_sc_hd__dfxtp_1
X_4225_ _5196_/Q input7/X _4234_/S vssd1 vssd1 vccd1 vccd1 _4226_/B sky130_fd_sc_hd__mux2_1
X_4156_ _5207_/Q _3531_/A _3665_/A vssd1 vssd1 vccd1 vccd1 _4156_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3107_ _5381_/Q _3028_/X _4834_/A _3009_/X _3106_/X vssd1 vssd1 vccd1 vccd1 _5381_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4087_ _4094_/A vssd1 vssd1 vccd1 vccd1 _4954_/A sky130_fd_sc_hd__buf_4
X_3038_ _3013_/B _3067_/B _3021_/A vssd1 vssd1 vccd1 vccd1 _3038_/X sky130_fd_sc_hd__o21a_1
XFILLER_36_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4989_ _5335_/CLK _4989_/D vssd1 vssd1 vccd1 vccd1 _4989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_3_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput15 io_in[30] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_2
Xinput26 la1_data_in[16] vssd1 vssd1 vccd1 vccd1 _5343_/D sky130_fd_sc_hd__clkbuf_1
Xinput37 la1_data_in[26] vssd1 vssd1 vccd1 vccd1 _5353_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4010_ _2743_/A _3705_/B _2736_/B vssd1 vssd1 vccd1 vccd1 _4010_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4912_ _5422_/Q _2902_/X _4916_/S vssd1 vssd1 vccd1 vccd1 _4913_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4843_ _5372_/D _4840_/X _4841_/Y _4842_/X vssd1 vssd1 vccd1 vccd1 _5404_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4774_ _5365_/Q _5364_/Q _4774_/C vssd1 vssd1 vccd1 vccd1 _4780_/C sky130_fd_sc_hd__and3_1
X_3725_ _3720_/X _3724_/Y _5019_/Q _3711_/X vssd1 vssd1 vccd1 vccd1 _5019_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3656_ _4837_/B vssd1 vssd1 vccd1 vccd1 _3656_/Y sky130_fd_sc_hd__inv_2
X_2607_ _2609_/A vssd1 vssd1 vccd1 vccd1 _2607_/Y sky130_fd_sc_hd__inv_2
X_3587_ _3673_/B _3662_/C vssd1 vssd1 vccd1 vccd1 _4434_/C sky130_fd_sc_hd__nor2_2
X_5326_ _5328_/CLK _5326_/D vssd1 vssd1 vccd1 vccd1 _5326_/Q sky130_fd_sc_hd__dfxtp_1
X_2538_ _2743_/A _2562_/A vssd1 vssd1 vccd1 vccd1 _2558_/A sky130_fd_sc_hd__and2_1
X_5257_ _5435_/CLK _5257_/D vssd1 vssd1 vccd1 vccd1 _5257_/Q sky130_fd_sc_hd__dfxtp_1
X_4208_ _4207_/X _5191_/Q _4214_/S vssd1 vssd1 vccd1 vccd1 _4209_/A sky130_fd_sc_hd__mux2_1
X_5188_ _5444_/CLK _5188_/D vssd1 vssd1 vccd1 vccd1 _5188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4139_ _4261_/S vssd1 vssd1 vccd1 vccd1 _4148_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_43_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5532__122 vssd1 vssd1 vccd1 vccd1 _5532__122/HI _5532__122/LO sky130_fd_sc_hd__conb_1
XFILLER_52_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3510_ _3510_/A _3510_/B _3510_/C vssd1 vssd1 vccd1 vccd1 _3526_/A sky130_fd_sc_hd__and3_1
X_4490_ _5265_/Q _5103_/Q _4492_/S vssd1 vssd1 vccd1 vccd1 _4491_/A sky130_fd_sc_hd__mux2_1
X_3441_ _3847_/A vssd1 vssd1 vccd1 vccd1 _3841_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3372_ _3372_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3373_/C sky130_fd_sc_hd__nor2_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5111_ _5111_/CLK _5111_/D vssd1 vssd1 vccd1 vccd1 _5111_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5245_/CLK _5042_/D vssd1 vssd1 vccd1 vccd1 _5042_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5516__106 vssd1 vssd1 vccd1 vccd1 _5516__106/HI _5632_/A sky130_fd_sc_hd__conb_1
XFILLER_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4826_ _4826_/A vssd1 vssd1 vccd1 vccd1 _5402_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4757_ _4757_/A _4757_/B vssd1 vssd1 vccd1 vccd1 _5359_/D sky130_fd_sc_hd__nor2_1
X_3708_ _3729_/B vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__clkbuf_2
X_4688_ _4692_/B _4692_/C vssd1 vssd1 vccd1 vccd1 _4694_/B sky130_fd_sc_hd__and2_1
X_3639_ _3639_/A vssd1 vssd1 vccd1 vccd1 _5001_/D sky130_fd_sc_hd__clkbuf_1
X_5309_ _5435_/CLK _5309_/D vssd1 vssd1 vccd1 vccd1 _5309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_21_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5371_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3990_ _5444_/Q vssd1 vssd1 vccd1 vccd1 _4203_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2941_ _3023_/A _2941_/B vssd1 vssd1 vccd1 vccd1 _4831_/B sky130_fd_sc_hd__xnor2_1
XFILLER_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2872_ _5030_/Q _5029_/Q _2872_/S vssd1 vssd1 vccd1 vccd1 _2872_/X sky130_fd_sc_hd__mux2_1
X_4611_ _4611_/A vssd1 vssd1 vccd1 vccd1 _4632_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5591_ _5591_/A _2621_/Y vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__ebufn_8
XFILLER_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4542_ _4542_/A vssd1 vssd1 vccd1 vccd1 _5284_/D sky130_fd_sc_hd__clkbuf_1
X_4473_ _5257_/Q hold144/X _4481_/S vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__mux2_1
X_3424_ _3424_/A _3442_/A _3424_/C vssd1 vssd1 vccd1 vccd1 _3749_/B sky130_fd_sc_hd__and3_1
X_3355_ _3355_/A _3355_/B vssd1 vssd1 vccd1 vccd1 _3356_/B sky130_fd_sc_hd__nor2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3442_/A _3772_/B _3286_/C vssd1 vssd1 vccd1 vccd1 _3409_/A sky130_fd_sc_hd__and3_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5058_/CLK _5025_/D vssd1 vssd1 vccd1 vccd1 _5025_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4809_ _4809_/A vssd1 vssd1 vccd1 vccd1 _5394_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3140_ _3074_/X _5384_/Q _3076_/X _5315_/Q vssd1 vssd1 vccd1 vccd1 _3141_/B sky130_fd_sc_hd__a22o_1
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3071_ _3139_/A _3071_/B vssd1 vssd1 vccd1 vccd1 _3083_/A sky130_fd_sc_hd__xnor2_1
X_3973_ _3980_/A vssd1 vssd1 vccd1 vccd1 _3973_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2924_ _2924_/A _5233_/Q vssd1 vssd1 vccd1 vccd1 _3027_/A sky130_fd_sc_hd__or2_1
X_2855_ _5022_/Q _5021_/Q _2859_/S vssd1 vssd1 vccd1 vccd1 _2855_/X sky130_fd_sc_hd__mux2_1
X_5574_ _5574_/A _2600_/Y vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__ebufn_8
X_4525_ _4525_/A vssd1 vssd1 vccd1 vccd1 _5276_/D sky130_fd_sc_hd__clkbuf_1
X_2786_ _5444_/Q _4508_/A _2786_/C _2786_/D vssd1 vssd1 vccd1 vccd1 _2787_/B sky130_fd_sc_hd__or4_2
X_4456_ _4450_/Y _4455_/X _4445_/X vssd1 vssd1 vccd1 vccd1 _4457_/C sky130_fd_sc_hd__o21ai_1
X_3407_ _3847_/A _3835_/A _3403_/X _3238_/A _3406_/Y vssd1 vssd1 vccd1 vccd1 _3408_/B
+ sky130_fd_sc_hd__a311o_1
X_4387_ _4400_/A _4387_/B vssd1 vssd1 vccd1 vccd1 _4387_/X sky130_fd_sc_hd__or2_1
X_3338_ _3338_/A vssd1 vssd1 vccd1 vccd1 _3343_/A sky130_fd_sc_hd__inv_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3269_ _3379_/A vssd1 vssd1 vccd1 vccd1 _3352_/S sky130_fd_sc_hd__dlymetal6s2s_1
X_5008_ _5444_/CLK _5008_/D vssd1 vssd1 vccd1 vccd1 _5008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2640_ _2640_/A vssd1 vssd1 vccd1 vccd1 _2640_/Y sky130_fd_sc_hd__inv_2
X_2571_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2571_/Y sky130_fd_sc_hd__inv_2
X_4310_ _4310_/A vssd1 vssd1 vccd1 vccd1 _5218_/D sky130_fd_sc_hd__clkbuf_1
X_5290_ _5437_/CLK _5290_/D vssd1 vssd1 vccd1 vccd1 _5290_/Q sky130_fd_sc_hd__dfxtp_1
X_4241_ _4241_/A vssd1 vssd1 vccd1 vccd1 _5200_/D sky130_fd_sc_hd__clkbuf_1
X_4172_ _4172_/A vssd1 vssd1 vccd1 vccd1 _5180_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3123_ _3187_/A _3648_/A vssd1 vssd1 vccd1 vccd1 _3123_/X sky130_fd_sc_hd__or2_1
XFILLER_27_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3054_ _3155_/B _5379_/Q _3053_/X _3129_/A vssd1 vssd1 vccd1 vccd1 _3055_/B sky130_fd_sc_hd__o211a_1
XFILLER_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3956_ _5091_/Q _3955_/X _3956_/S vssd1 vssd1 vccd1 vccd1 _3957_/A sky130_fd_sc_hd__mux2_1
X_2907_ _2953_/B _2907_/B _2977_/C vssd1 vssd1 vccd1 vccd1 _2907_/X sky130_fd_sc_hd__or3_1
X_5626_ _5629_/A _2663_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[22] sky130_fd_sc_hd__ebufn_8
X_3887_ _3887_/A vssd1 vssd1 vccd1 vccd1 _5076_/D sky130_fd_sc_hd__clkbuf_1
X_2838_ _2838_/A vssd1 vssd1 vccd1 vccd1 _2838_/X sky130_fd_sc_hd__clkbuf_2
X_5557_ _5557_/A _2581_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[23] sky130_fd_sc_hd__ebufn_8
X_2769_ _2769_/A vssd1 vssd1 vccd1 vccd1 _5148_/D sky130_fd_sc_hd__buf_2
X_4508_ _4508_/A _4508_/B _4508_/C vssd1 vssd1 vccd1 vccd1 _4514_/B sky130_fd_sc_hd__or3_2
X_4439_ _4450_/A _4438_/Y _2766_/A vssd1 vssd1 vccd1 vccd1 _4439_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_59_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3810_ _5048_/Q _5047_/Q _3810_/C vssd1 vssd1 vccd1 vccd1 _3813_/B sky130_fd_sc_hd__and3_1
X_4790_ _4790_/A vssd1 vssd1 vccd1 vccd1 _5370_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3741_ _3750_/A vssd1 vssd1 vccd1 vccd1 _3741_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_18 _5353_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_29 _2766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3672_ _3672_/A vssd1 vssd1 vccd1 vccd1 _5005_/D sky130_fd_sc_hd__clkbuf_1
X_2623_ _2635_/A vssd1 vssd1 vccd1 vccd1 _2628_/A sky130_fd_sc_hd__buf_4
X_5411_ _5403_/Q _5411_/D vssd1 vssd1 vccd1 vccd1 _5411_/Q sky130_fd_sc_hd__dfxtp_1
X_5342_ _5351_/CLK _5342_/D vssd1 vssd1 vccd1 vccd1 _5342_/Q sky130_fd_sc_hd__dfxtp_1
X_2554_ _2554_/A _2554_/B vssd1 vssd1 vccd1 vccd1 _5114_/D sky130_fd_sc_hd__nor2_1
X_5273_ _5322_/CLK _5273_/D vssd1 vssd1 vccd1 vccd1 _5273_/Q sky130_fd_sc_hd__dfxtp_1
X_4224_ _4224_/A vssd1 vssd1 vccd1 vccd1 _5195_/D sky130_fd_sc_hd__clkbuf_1
X_4155_ _5178_/Q _5179_/Q _5177_/Q vssd1 vssd1 vccd1 vccd1 _4155_/X sky130_fd_sc_hd__or3b_2
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3106_ _3106_/A _5237_/Q vssd1 vssd1 vccd1 vccd1 _3106_/X sky130_fd_sc_hd__or2_1
X_4086_ _4086_/A _4086_/B vssd1 vssd1 vccd1 vccd1 _5152_/D sky130_fd_sc_hd__nor2_1
X_3037_ _3066_/B vssd1 vssd1 vccd1 vccd1 _3040_/A sky130_fd_sc_hd__inv_2
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4988_ _5335_/CLK _4988_/D vssd1 vssd1 vccd1 vccd1 _4988_/Q sky130_fd_sc_hd__dfxtp_1
X_3939_ _5262_/Q _3915_/A _3699_/A _5288_/Q vssd1 vssd1 vccd1 vccd1 _3939_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5609_ _5609_/A _2643_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[5] sky130_fd_sc_hd__ebufn_8
XFILLER_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput27 la1_data_in[17] vssd1 vssd1 vccd1 vccd1 _5344_/D sky130_fd_sc_hd__clkbuf_1
Xinput16 io_in[31] vssd1 vssd1 vccd1 vccd1 _4978_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput38 la1_data_in[28] vssd1 vssd1 vccd1 vccd1 _2786_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_38_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4911_ _4911_/A vssd1 vssd1 vccd1 vccd1 _5421_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_18_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4842_ _4902_/A vssd1 vssd1 vccd1 vccd1 _4842_/X sky130_fd_sc_hd__clkbuf_2
X_4773_ _4773_/A _4773_/B vssd1 vssd1 vccd1 vccd1 _5364_/D sky130_fd_sc_hd__nor2_1
X_3724_ _3724_/A _3724_/B vssd1 vssd1 vccd1 vccd1 _3724_/Y sky130_fd_sc_hd__nand2_1
X_3655_ _3655_/A _3655_/B vssd1 vssd1 vccd1 vccd1 _4837_/B sky130_fd_sc_hd__xnor2_4
X_2606_ _2609_/A vssd1 vssd1 vccd1 vccd1 _2606_/Y sky130_fd_sc_hd__inv_2
X_3586_ _3592_/A _3510_/C _3682_/C vssd1 vssd1 vccd1 vccd1 _3586_/Y sky130_fd_sc_hd__o21ai_1
X_5325_ _5328_/CLK _5325_/D vssd1 vssd1 vccd1 vccd1 _5325_/Q sky130_fd_sc_hd__dfxtp_1
X_2537_ _3705_/B _5110_/Q _2560_/B vssd1 vssd1 vccd1 vccd1 _2562_/A sky130_fd_sc_hd__and3_1
X_5256_ _5305_/CLK _5256_/D vssd1 vssd1 vccd1 vccd1 _5256_/Q sky130_fd_sc_hd__dfxtp_1
X_4207_ _5415_/Q _5366_/Q _4216_/S vssd1 vssd1 vccd1 vccd1 _4207_/X sky130_fd_sc_hd__mux2_1
XFILLER_56_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5187_ _5444_/CLK _5187_/D vssd1 vssd1 vccd1 vccd1 _5187_/Q sky130_fd_sc_hd__dfxtp_1
X_4138_ _4138_/A vssd1 vssd1 vccd1 vccd1 _5170_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_28_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4069_ _5383_/Q hold67/A _4071_/S vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_137_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3440_ _3440_/A vssd1 vssd1 vccd1 vccd1 _5594_/A sky130_fd_sc_hd__clkbuf_1
X_3371_ _3379_/A vssd1 vssd1 vccd1 vccd1 _3374_/A sky130_fd_sc_hd__inv_2
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5110_ _5110_/CLK _5110_/D vssd1 vssd1 vccd1 vccd1 _5110_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5245_/CLK _5041_/D vssd1 vssd1 vccd1 vccd1 _5041_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
XFILLER_53_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4825_ _4837_/B _5402_/Q _4825_/S vssd1 vssd1 vccd1 vccd1 _4826_/A sky130_fd_sc_hd__mux2_1
X_4756_ _5359_/Q _4758_/C _4746_/X vssd1 vssd1 vccd1 vccd1 _4757_/B sky130_fd_sc_hd__o21ai_1
X_3707_ _3726_/A _3726_/B _3707_/C_N vssd1 vssd1 vccd1 vccd1 _3707_/X sky130_fd_sc_hd__or3b_1
X_4687_ _3894_/B _4680_/X _4681_/X _4553_/A _4093_/A vssd1 vssd1 vccd1 vccd1 _5323_/D
+ sky130_fd_sc_hd__a221o_1
X_3638_ _3637_/X _3891_/B _3643_/S vssd1 vssd1 vccd1 vccd1 _3639_/A sky130_fd_sc_hd__mux2_1
X_3569_ _3569_/A vssd1 vssd1 vccd1 vccd1 _3569_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5308_ _5435_/CLK _5308_/D vssd1 vssd1 vccd1 vccd1 _5308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5487__77 vssd1 vssd1 vccd1 vccd1 _5487__77/HI _5565_/A sky130_fd_sc_hd__conb_1
X_5239_ _5445_/CLK _5239_/D vssd1 vssd1 vccd1 vccd1 _5239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_12_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2940_ _2938_/A _2939_/Y _2994_/A vssd1 vssd1 vccd1 vccd1 _2941_/B sky130_fd_sc_hd__mux2_1
X_2871_ _3476_/A _2868_/X _2869_/X _3476_/B _4034_/B vssd1 vssd1 vccd1 vccd1 _2871_/X
+ sky130_fd_sc_hd__a221o_1
X_4610_ _4610_/A vssd1 vssd1 vccd1 vccd1 _5305_/D sky130_fd_sc_hd__clkbuf_1
X_5590_ _5590_/A _2620_/Y vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__ebufn_8
X_4541_ _5284_/Q _5431_/Q _4541_/S vssd1 vssd1 vccd1 vccd1 _4542_/A sky130_fd_sc_hd__mux2_1
X_4472_ _4549_/S vssd1 vssd1 vccd1 vccd1 _4481_/S sky130_fd_sc_hd__clkbuf_2
X_3423_ _3853_/A _3851_/A vssd1 vssd1 vccd1 vccd1 _3427_/A sky130_fd_sc_hd__or2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3354_/A _3354_/B vssd1 vssd1 vccd1 vccd1 _3355_/A sky130_fd_sc_hd__nor2_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3285_ _3424_/C _3285_/B vssd1 vssd1 vccd1 vccd1 _3286_/C sky130_fd_sc_hd__or2_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5032_/CLK _5024_/D vssd1 vssd1 vccd1 vccd1 _5024_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4808_ _4832_/C _5394_/Q _4812_/S vssd1 vssd1 vccd1 vccd1 _4809_/A sky130_fd_sc_hd__mux2_1
X_4739_ _4739_/A _4739_/B vssd1 vssd1 vccd1 vccd1 _5354_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3070_ _3108_/A _5395_/Q vssd1 vssd1 vccd1 vccd1 _3071_/B sky130_fd_sc_hd__and2_1
XFILLER_48_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3972_ _4906_/A vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2923_ _5243_/Q vssd1 vssd1 vccd1 vccd1 _2924_/A sky130_fd_sc_hd__inv_2
XFILLER_31_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2854_ _4034_/B vssd1 vssd1 vccd1 vccd1 _2854_/Y sky130_fd_sc_hd__inv_2
X_2785_ _2785_/A _2785_/B _2785_/C _2785_/D vssd1 vssd1 vccd1 vccd1 _2790_/B sky130_fd_sc_hd__or4_2
X_5573_ _5573_/A _2599_/Y vssd1 vssd1 vccd1 vccd1 io_out[7] sky130_fd_sc_hd__ebufn_8
X_4524_ _5276_/Q _5423_/Q _4530_/S vssd1 vssd1 vccd1 vccd1 _4525_/A sky130_fd_sc_hd__mux2_1
X_4455_ _5252_/Q _4455_/B vssd1 vssd1 vccd1 vccd1 _4455_/X sky130_fd_sc_hd__and2_1
X_3406_ _3824_/B _3824_/C vssd1 vssd1 vccd1 vccd1 _3406_/Y sky130_fd_sc_hd__nand2_1
X_4386_ _5196_/Q _5166_/Q _4399_/S vssd1 vssd1 vccd1 vccd1 _4387_/B sky130_fd_sc_hd__mux2_1
X_3337_ _3337_/A _3337_/B vssd1 vssd1 vccd1 vccd1 _3338_/A sky130_fd_sc_hd__or2_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5457__47 vssd1 vssd1 vccd1 vccd1 _5457__47/HI _5534_/A sky130_fd_sc_hd__conb_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _3268_/A _3337_/A vssd1 vssd1 vccd1 vccd1 _3379_/A sky130_fd_sc_hd__xor2_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3199_ _5054_/Q vssd1 vssd1 vccd1 vccd1 _3823_/B sky130_fd_sc_hd__inv_2
X_5007_ _5369_/CLK _5007_/D vssd1 vssd1 vccd1 vccd1 _5007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5471__61 vssd1 vssd1 vccd1 vccd1 _5471__61/HI _5548_/A sky130_fd_sc_hd__conb_1
XFILLER_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2570_ _2572_/A vssd1 vssd1 vccd1 vccd1 _2570_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4240_ _4252_/A _4240_/B vssd1 vssd1 vccd1 vccd1 _4241_/A sky130_fd_sc_hd__and2_1
X_4171_ _4170_/X _5180_/Q _4180_/S vssd1 vssd1 vccd1 vccd1 _4172_/A sky130_fd_sc_hd__mux2_1
X_3122_ _3139_/A vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__clkbuf_4
X_3053_ _5310_/Q _3075_/B _2952_/Y input45/X _3074_/A vssd1 vssd1 vccd1 vccd1 _3053_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3955_ _5265_/Q _3915_/A _3943_/X _5087_/Q _3947_/X vssd1 vssd1 vccd1 vccd1 _3955_/X
+ sky130_fd_sc_hd__a221o_1
X_2906_ _2906_/A _2906_/B _2906_/C _2906_/D vssd1 vssd1 vccd1 vccd1 _2977_/C sky130_fd_sc_hd__or4_1
X_5625_ _5625_/A _2662_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[21] sky130_fd_sc_hd__ebufn_8
X_3886_ hold4/A _3186_/X _3888_/S vssd1 vssd1 vccd1 vccd1 _3887_/A sky130_fd_sc_hd__mux2_1
X_2837_ _2832_/X _2836_/Y _2843_/S vssd1 vssd1 vccd1 vccd1 _2837_/X sky130_fd_sc_hd__a21o_1
X_5556_ _5556_/A _2578_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[22] sky130_fd_sc_hd__ebufn_8
X_2768_ _2768_/A _2768_/B vssd1 vssd1 vccd1 vccd1 _2769_/A sky130_fd_sc_hd__and2_1
X_4507_ _5301_/Q _3913_/A _4506_/Y _3912_/B vssd1 vssd1 vccd1 vccd1 _4508_/C sky130_fd_sc_hd__a22o_1
X_2699_ _4508_/A vssd1 vssd1 vccd1 vccd1 _4115_/A sky130_fd_sc_hd__buf_2
X_4438_ _4438_/A _4438_/B vssd1 vssd1 vccd1 vccd1 _4438_/Y sky130_fd_sc_hd__nor2_1
X_4369_ input7/X _5162_/Q _4380_/S vssd1 vssd1 vccd1 vccd1 _4370_/B sky130_fd_sc_hd__mux2_1
XFILLER_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3740_ _3740_/A vssd1 vssd1 vccd1 vccd1 _3740_/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_19 _5582_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3671_ _3670_/X _5005_/Q _3675_/S vssd1 vssd1 vccd1 vccd1 _3672_/A sky130_fd_sc_hd__mux2_1
X_5410_ _5403_/Q _5410_/D vssd1 vssd1 vccd1 vccd1 _5410_/Q sky130_fd_sc_hd__dfxtp_1
X_2622_ _2622_/A vssd1 vssd1 vccd1 vccd1 _2622_/Y sky130_fd_sc_hd__inv_2
X_5341_ _5351_/CLK _5341_/D vssd1 vssd1 vccd1 vccd1 _5341_/Q sky130_fd_sc_hd__dfxtp_1
X_2553_ _5114_/Q _2556_/A _2544_/X vssd1 vssd1 vccd1 vccd1 _2554_/B sky130_fd_sc_hd__o21ai_1
X_5272_ _5323_/CLK _5272_/D vssd1 vssd1 vccd1 vccd1 _5272_/Q sky130_fd_sc_hd__dfxtp_1
X_4223_ _4235_/A _4223_/B vssd1 vssd1 vccd1 vccd1 _4224_/A sky130_fd_sc_hd__and2_1
X_4154_ _4154_/A vssd1 vssd1 vccd1 vccd1 _4421_/S sky130_fd_sc_hd__clkbuf_2
X_4085_ _5152_/Q _4083_/A _4081_/X vssd1 vssd1 vccd1 vccd1 _4086_/B sky130_fd_sc_hd__o21ai_1
X_3105_ _3154_/A _3105_/B vssd1 vssd1 vccd1 vccd1 _4834_/A sky130_fd_sc_hd__xnor2_4
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3036_ _3036_/A _3036_/B vssd1 vssd1 vccd1 vccd1 _3066_/B sky130_fd_sc_hd__and2_1
XFILLER_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4987_ _5335_/CLK _4987_/D vssd1 vssd1 vccd1 vccd1 _4987_/Q sky130_fd_sc_hd__dfxtp_1
X_3938_ _5087_/Q _3932_/X _3937_/X vssd1 vssd1 vccd1 vccd1 _5087_/D sky130_fd_sc_hd__o21a_1
XFILLER_137_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3869_ hold31/A _4833_/A _3873_/S vssd1 vssd1 vccd1 vccd1 _3870_/A sky130_fd_sc_hd__mux2_1
X_5608_ _5608_/A _2640_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[4] sky130_fd_sc_hd__ebufn_8
XFILLER_11_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5539_ _5539_/A _2688_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[5] sky130_fd_sc_hd__ebufn_8
Xclkbuf_leaf_15_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5436_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_59_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput28 la1_data_in[18] vssd1 vssd1 vccd1 vccd1 _5345_/D sky130_fd_sc_hd__clkbuf_1
Xinput17 io_in[32] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
Xinput39 la1_data_in[2] vssd1 vssd1 vccd1 vccd1 _2929_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4910_ _5421_/Q _2977_/A _4916_/S vssd1 vssd1 vccd1 vccd1 _4911_/A sky130_fd_sc_hd__mux2_1
XFILLER_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4841_ _5404_/Q _4841_/B vssd1 vssd1 vccd1 vccd1 _4841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4772_ _5364_/Q _4774_/C _4762_/X vssd1 vssd1 vccd1 vccd1 _4773_/B sky130_fd_sc_hd__o21ai_1
X_3723_ _3720_/X _3722_/Y _5018_/Q _3711_/X vssd1 vssd1 vccd1 vccd1 _5018_/D sky130_fd_sc_hd__o2bb2a_1
XFILLER_9_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3654_ _3654_/A _3654_/B vssd1 vssd1 vccd1 vccd1 _3655_/B sky130_fd_sc_hd__xnor2_2
X_2605_ _2609_/A vssd1 vssd1 vccd1 vccd1 _2605_/Y sky130_fd_sc_hd__inv_2
X_3585_ _4996_/Q _3583_/A _3584_/Y vssd1 vssd1 vccd1 vccd1 _4996_/D sky130_fd_sc_hd__o21a_1
X_5324_ _5328_/CLK _5324_/D vssd1 vssd1 vccd1 vccd1 _5324_/Q sky130_fd_sc_hd__dfxtp_1
X_2536_ _5111_/Q vssd1 vssd1 vccd1 vccd1 _3705_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5255_ _5305_/CLK _5255_/D vssd1 vssd1 vccd1 vccd1 _5255_/Q sky130_fd_sc_hd__dfxtp_1
X_4206_ _4206_/A vssd1 vssd1 vccd1 vccd1 _5190_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5186_ _5444_/CLK _5186_/D vssd1 vssd1 vccd1 vccd1 _5186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4137_ _5347_/Q _5170_/Q _4137_/S vssd1 vssd1 vccd1 vccd1 _4138_/A sky130_fd_sc_hd__mux2_1
XFILLER_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4068_ _4068_/A vssd1 vssd1 vccd1 vccd1 _5145_/D sky130_fd_sc_hd__clkbuf_1
X_3019_ _3020_/A _3020_/B vssd1 vssd1 vccd1 vccd1 _3021_/A sky130_fd_sc_hd__or2_1
XFILLER_24_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3370_ _3379_/A _3374_/B _3267_/X vssd1 vssd1 vccd1 vccd1 _3370_/X sky130_fd_sc_hd__o21ba_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5439_/CLK _5040_/D vssd1 vssd1 vccd1 vccd1 _5040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4824_ _4824_/A vssd1 vssd1 vccd1 vccd1 _5401_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4755_ _5359_/Q _4758_/C vssd1 vssd1 vccd1 vccd1 _4757_/A sky130_fd_sc_hd__and2_1
X_3706_ _3709_/A vssd1 vssd1 vccd1 vccd1 _3726_/B sky130_fd_sc_hd__clkbuf_2
X_4686_ _4686_/A vssd1 vssd1 vccd1 vccd1 _5322_/D sky130_fd_sc_hd__clkbuf_1
X_3637_ _3912_/B _3627_/X _3892_/B _3699_/A _3636_/Y vssd1 vssd1 vccd1 vccd1 _3637_/X
+ sky130_fd_sc_hd__a311o_1
X_3568_ _3572_/A _3575_/B vssd1 vssd1 vccd1 vccd1 _3571_/A sky130_fd_sc_hd__and2_1
XFILLER_0_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5307_ _5435_/CLK _5307_/D vssd1 vssd1 vccd1 vccd1 _5307_/Q sky130_fd_sc_hd__dfxtp_1
X_2519_ _5041_/Q vssd1 vssd1 vccd1 vccd1 _3788_/A sky130_fd_sc_hd__inv_2
X_3499_ _5246_/Q vssd1 vssd1 vccd1 vccd1 _3662_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5238_ _5436_/CLK _5238_/D vssd1 vssd1 vccd1 vccd1 _5238_/Q sky130_fd_sc_hd__dfxtp_2
X_5169_ _5351_/CLK _5169_/D vssd1 vssd1 vccd1 vccd1 _5169_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_29_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _4000_/A
+ sky130_fd_sc_hd__clkbuf_16
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_58_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2870_ _2870_/A _2870_/B vssd1 vssd1 vccd1 vccd1 _3476_/B sky130_fd_sc_hd__nor2_2
XFILLER_30_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4540_ _4540_/A vssd1 vssd1 vccd1 vccd1 _5283_/D sky130_fd_sc_hd__clkbuf_1
X_4471_ _4471_/A vssd1 vssd1 vccd1 vccd1 _4549_/S sky130_fd_sc_hd__clkbuf_2
X_3422_ _5060_/Q vssd1 vssd1 vccd1 vccd1 _3851_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5522__112 vssd1 vssd1 vccd1 vccd1 _5522__112/HI _5638_/A sky130_fd_sc_hd__conb_1
X_3353_ _3267_/X _3340_/Y _3352_/X vssd1 vssd1 vccd1 vccd1 _3353_/X sky130_fd_sc_hd__o21ba_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3284_/A vssd1 vssd1 vccd1 vccd1 _3772_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5058_/CLK _5023_/D vssd1 vssd1 vccd1 vccd1 _5023_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4807_ _4807_/A vssd1 vssd1 vccd1 vccd1 _5393_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_22_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2999_ _3033_/A _2999_/B vssd1 vssd1 vccd1 vccd1 _3002_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4738_ _4954_/A _4738_/B _5371_/D vssd1 vssd1 vccd1 vccd1 _5337_/D sky130_fd_sc_hd__nor3_1
X_4669_ _4587_/A _4328_/A _4589_/A _4586_/X _3691_/Y vssd1 vssd1 vccd1 vccd1 _4669_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3971_ _5095_/Q _3966_/X _5437_/D _2965_/X vssd1 vssd1 vccd1 vccd1 _5095_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2922_ _2922_/A vssd1 vssd1 vccd1 vccd1 _5372_/D sky130_fd_sc_hd__clkbuf_1
X_5641_ _5641_/A _2681_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[37] sky130_fd_sc_hd__ebufn_8
X_2853_ _5130_/Q vssd1 vssd1 vccd1 vccd1 _4034_/B sky130_fd_sc_hd__buf_2
X_5572_ _5572_/A _2597_/Y vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__ebufn_8
X_2784_ _4084_/B _2778_/A _2783_/Y _2717_/X _2720_/C vssd1 vssd1 vccd1 vccd1 _2785_/D
+ sky130_fd_sc_hd__a221o_1
X_4523_ _4523_/A vssd1 vssd1 vccd1 vccd1 _5275_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_7_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4454_ _4450_/A _4450_/B _4455_/B _5252_/Q vssd1 vssd1 vccd1 vccd1 _4457_/B sky130_fd_sc_hd__a31o_1
X_3405_ _3424_/A vssd1 vssd1 vccd1 vccd1 _3824_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_4385_ _4421_/S vssd1 vssd1 vccd1 vccd1 _4399_/S sky130_fd_sc_hd__clkbuf_2
X_3336_ _3336_/A _3349_/A vssd1 vssd1 vccd1 vccd1 _3337_/B sky130_fd_sc_hd__and2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3267_/A vssd1 vssd1 vccd1 vccd1 _3267_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5006_ _5245_/CLK _5006_/D vssd1 vssd1 vccd1 vccd1 _5006_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3198_ _5055_/Q vssd1 vssd1 vccd1 vccd1 _3823_/A sky130_fd_sc_hd__inv_2
XFILLER_14_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4170_ _5404_/Q _5355_/Q _4182_/S vssd1 vssd1 vccd1 vccd1 _4170_/X sky130_fd_sc_hd__mux2_1
X_3121_ _4791_/A vssd1 vssd1 vccd1 vccd1 _3187_/A sky130_fd_sc_hd__clkbuf_1
X_3052_ _3126_/A _5394_/Q _3126_/B vssd1 vssd1 vccd1 vccd1 _3057_/B sky130_fd_sc_hd__a21oi_1
XFILLER_36_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3954_ _5090_/Q _3932_/X _3953_/X _3642_/B vssd1 vssd1 vccd1 vccd1 _5090_/D sky130_fd_sc_hd__o22a_1
X_3885_ _3885_/A vssd1 vssd1 vccd1 vccd1 _5075_/D sky130_fd_sc_hd__clkbuf_1
X_2905_ _5600_/A _4964_/A _2953_/C vssd1 vssd1 vccd1 vccd1 _2905_/X sky130_fd_sc_hd__a21o_1
X_2836_ _3466_/A _2835_/Y _2817_/S vssd1 vssd1 vccd1 vccd1 _2836_/Y sky130_fd_sc_hd__a21oi_1
X_5624_ _5624_/A _2661_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[20] sky130_fd_sc_hd__ebufn_8
X_2767_ _2767_/A vssd1 vssd1 vccd1 vccd1 _5037_/D sky130_fd_sc_hd__clkbuf_1
X_5555_ _5555_/A _2577_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[21] sky130_fd_sc_hd__ebufn_8
X_2698_ _2698_/A vssd1 vssd1 vccd1 vccd1 _2698_/Y sky130_fd_sc_hd__inv_2
X_4506_ _4551_/B _4506_/B vssd1 vssd1 vccd1 vccd1 _4506_/Y sky130_fd_sc_hd__nand2_2
X_4437_ _4437_/A vssd1 vssd1 vccd1 vccd1 _4438_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _5228_/Q _4362_/X _4367_/X _2750_/X vssd1 vssd1 vccd1 vccd1 _5228_/D sky130_fd_sc_hd__o211a_1
X_3319_ _3319_/A _3319_/B _3319_/C vssd1 vssd1 vccd1 vccd1 _3321_/A sky130_fd_sc_hd__and3_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _5166_/Q _4285_/X _4276_/A _5192_/Q vssd1 vssd1 vccd1 vccd1 _4299_/X sky130_fd_sc_hd__a22o_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3670_ _3533_/A _4165_/A _3667_/B _3682_/D _3669_/Y vssd1 vssd1 vccd1 vccd1 _3670_/X
+ sky130_fd_sc_hd__a311o_1
X_2621_ _2622_/A vssd1 vssd1 vccd1 vccd1 _2621_/Y sky130_fd_sc_hd__inv_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5340_ _5351_/CLK _5340_/D vssd1 vssd1 vccd1 vccd1 _5340_/Q sky130_fd_sc_hd__dfxtp_1
X_2552_ _2736_/B _2743_/A _2562_/A vssd1 vssd1 vccd1 vccd1 _2556_/A sky130_fd_sc_hd__and3_1
X_5271_ _5323_/CLK _5271_/D vssd1 vssd1 vccd1 vccd1 _5271_/Q sky130_fd_sc_hd__dfxtp_1
X_4222_ _5195_/Q input6/X _4234_/S vssd1 vssd1 vccd1 vccd1 _4223_/B sky130_fd_sc_hd__mux2_1
X_4153_ _5248_/Q _4730_/B vssd1 vssd1 vccd1 vccd1 _4154_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4084_ _5152_/Q _4084_/B _4092_/B vssd1 vssd1 vccd1 vccd1 _4086_/A sky130_fd_sc_hd__and3_1
X_3104_ _3646_/A _3101_/Y _3102_/X _3103_/X vssd1 vssd1 vccd1 vccd1 _3105_/B sky130_fd_sc_hd__o31a_2
X_3035_ _3035_/A _3035_/B vssd1 vssd1 vccd1 vccd1 _3036_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4986_ _5446_/CLK _4986_/D vssd1 vssd1 vccd1 vccd1 _5585_/A sky130_fd_sc_hd__dfxtp_4
X_3937_ _5287_/Q _3910_/X _3697_/A _3936_/X vssd1 vssd1 vccd1 vccd1 _3937_/X sky130_fd_sc_hd__a211o_1
XFILLER_32_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3868_ _3868_/A vssd1 vssd1 vccd1 vccd1 _5067_/D sky130_fd_sc_hd__clkbuf_1
X_5607_ _5607_/A _2639_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[3] sky130_fd_sc_hd__ebufn_8
X_3799_ _3799_/A vssd1 vssd1 vccd1 vccd1 _5044_/D sky130_fd_sc_hd__clkbuf_1
X_2819_ _5131_/Q _2822_/B vssd1 vssd1 vccd1 vccd1 _2827_/C sky130_fd_sc_hd__or2_1
XFILLER_11_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5538_ _5538_/A _2687_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[4] sky130_fd_sc_hd__ebufn_8
XFILLER_47_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 io_in[33] vssd1 vssd1 vccd1 vccd1 _4982_/A sky130_fd_sc_hd__clkbuf_2
Xinput29 la1_data_in[19] vssd1 vssd1 vccd1 vccd1 _5346_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_2_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4840_ _4841_/B vssd1 vssd1 vccd1 vccd1 _4840_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4771_ _5364_/Q _5363_/Q _4771_/C vssd1 vssd1 vccd1 vccd1 _4773_/A sky130_fd_sc_hd__and3_1
X_3722_ _3722_/A _3724_/B vssd1 vssd1 vccd1 vccd1 _3722_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3653_ _3649_/B _3649_/Y _3653_/S vssd1 vssd1 vccd1 vccd1 _3654_/B sky130_fd_sc_hd__mux2_1
X_2604_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2609_/A sky130_fd_sc_hd__clkbuf_2
X_3584_ _4996_/Q _3583_/A _3569_/A vssd1 vssd1 vccd1 vccd1 _3584_/Y sky130_fd_sc_hd__a21boi_1
X_5323_ _5323_/CLK _5323_/D vssd1 vssd1 vccd1 vccd1 _5323_/Q sky130_fd_sc_hd__dfxtp_1
X_2535_ _5112_/Q vssd1 vssd1 vccd1 vccd1 _2743_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5254_ _5322_/CLK _5254_/D vssd1 vssd1 vccd1 vccd1 _5254_/Q sky130_fd_sc_hd__dfxtp_1
X_5185_ _5444_/CLK _5185_/D vssd1 vssd1 vccd1 vccd1 _5185_/Q sky130_fd_sc_hd__dfxtp_1
X_4205_ _4204_/X _5190_/Q _4214_/S vssd1 vssd1 vccd1 vccd1 _4206_/A sky130_fd_sc_hd__mux2_1
X_4136_ _4136_/A vssd1 vssd1 vccd1 vccd1 _5169_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4067_ _5382_/Q hold76/A _4071_/S vssd1 vssd1 vccd1 vccd1 _4068_/A sky130_fd_sc_hd__mux2_1
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3018_ _3130_/A _3018_/B vssd1 vssd1 vccd1 vccd1 _3020_/B sky130_fd_sc_hd__xnor2_1
XFILLER_24_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4969_ _2942_/X _4965_/Y _4968_/X _4902_/X vssd1 vssd1 vccd1 vccd1 _5448_/D sky130_fd_sc_hd__o211a_1
XFILLER_137_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5501__91 vssd1 vssd1 vccd1 vccd1 _5501__91/HI _5604_/A sky130_fd_sc_hd__conb_1
XFILLER_19_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_0_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5245_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4823_ _3186_/X _5401_/Q _4823_/S vssd1 vssd1 vccd1 vccd1 _4824_/A sky130_fd_sc_hd__mux2_1
X_4754_ _4758_/C _4754_/B vssd1 vssd1 vccd1 vccd1 _5358_/D sky130_fd_sc_hd__nor2_1
X_3705_ _3705_/A _3705_/B _3705_/C _3705_/D vssd1 vssd1 vccd1 vccd1 _3709_/A sky130_fd_sc_hd__nor4_1
X_4685_ _4685_/A _4685_/B vssd1 vssd1 vccd1 vccd1 _4686_/A sky130_fd_sc_hd__or2_1
X_3636_ _3642_/A _3891_/B vssd1 vssd1 vccd1 vccd1 _3636_/Y sky130_fd_sc_hd__xnor2_1
X_3567_ _3567_/A vssd1 vssd1 vccd1 vccd1 _4990_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2518_ _5042_/Q _5041_/Q vssd1 vssd1 vccd1 vccd1 _2518_/Y sky130_fd_sc_hd__xnor2_1
X_5306_ _5436_/CLK _5306_/D vssd1 vssd1 vccd1 vccd1 _5306_/Q sky130_fd_sc_hd__dfxtp_1
X_3498_ _3498_/A vssd1 vssd1 vccd1 vccd1 _5575_/A sky130_fd_sc_hd__clkbuf_1
X_5237_ _5445_/CLK _5237_/D vssd1 vssd1 vccd1 vccd1 _5237_/Q sky130_fd_sc_hd__dfxtp_1
X_5168_ _5351_/CLK _5168_/D vssd1 vssd1 vccd1 vccd1 _5168_/Q sky130_fd_sc_hd__dfxtp_1
X_4119_ _4119_/A vssd1 vssd1 vccd1 vccd1 _5161_/D sky130_fd_sc_hd__clkbuf_1
X_5099_ _5435_/CLK _5099_/D vssd1 vssd1 vccd1 vccd1 _5099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5478__68 vssd1 vssd1 vccd1 vccd1 _5478__68/HI _5555_/A sky130_fd_sc_hd__conb_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_59_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4470_ _4470_/A vssd1 vssd1 vccd1 vccd1 _5256_/D sky130_fd_sc_hd__clkbuf_1
X_3421_ _5061_/Q vssd1 vssd1 vccd1 vccd1 _3853_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3352_ _3374_/B _3351_/X _3352_/S vssd1 vssd1 vccd1 vccd1 _3352_/X sky130_fd_sc_hd__mux2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _5057_/Q vssd1 vssd1 vccd1 vccd1 _3442_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _5032_/CLK _5022_/D vssd1 vssd1 vccd1 vccd1 _5022_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5492__82 vssd1 vssd1 vccd1 vccd1 _5492__82/HI _5570_/A sky130_fd_sc_hd__conb_1
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4806_ _4833_/A _5393_/Q _4812_/S vssd1 vssd1 vccd1 vccd1 _4807_/A sky130_fd_sc_hd__mux2_1
XFILLER_22_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2998_ _5240_/Q _5376_/Q _2997_/X _2910_/A vssd1 vssd1 vccd1 vccd1 _2999_/B sky130_fd_sc_hd__o211a_1
X_4737_ _4737_/A vssd1 vssd1 vccd1 vccd1 _5371_/D sky130_fd_sc_hd__buf_2
X_4668_ _4668_/A vssd1 vssd1 vccd1 vccd1 _5318_/D sky130_fd_sc_hd__clkbuf_1
X_3619_ _5323_/Q _3893_/B vssd1 vssd1 vccd1 vccd1 _3912_/B sky130_fd_sc_hd__or2_2
XFILLER_1_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4599_ _4666_/S vssd1 vssd1 vccd1 vccd1 _4617_/S sky130_fd_sc_hd__buf_2
XFILLER_0_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3970_ _5094_/Q _3966_/X _5437_/D _2942_/X vssd1 vssd1 vccd1 vccd1 _5094_/D sky130_fd_sc_hd__a22o_1
XFILLER_23_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2921_ _5228_/Q _2919_/X _4791_/A vssd1 vssd1 vccd1 vccd1 _2922_/A sky130_fd_sc_hd__mux2_1
XFILLER_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _5640_/A _2680_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[36] sky130_fd_sc_hd__ebufn_8
X_2852_ _3489_/A _4042_/A vssd1 vssd1 vccd1 vccd1 _2852_/Y sky130_fd_sc_hd__nor2_1
X_5571_ _5571_/A _2596_/Y vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__ebufn_8
X_2783_ _5152_/Q _5151_/Q vssd1 vssd1 vccd1 vccd1 _2783_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4522_ _5275_/Q _5422_/Q _4530_/S vssd1 vssd1 vccd1 vccd1 _4523_/A sky130_fd_sc_hd__mux2_1
X_4453_ _4739_/B _4453_/B vssd1 vssd1 vccd1 vccd1 _5251_/D sky130_fd_sc_hd__nor2_1
X_3404_ _5059_/Q vssd1 vssd1 vccd1 vccd1 _3824_/B sky130_fd_sc_hd__clkbuf_1
X_4384_ _4422_/A vssd1 vssd1 vccd1 vccd1 _4400_/A sky130_fd_sc_hd__clkbuf_1
X_3335_ _3551_/B _3358_/A _3344_/A _3357_/A vssd1 vssd1 vccd1 vccd1 _3390_/B sky130_fd_sc_hd__or4_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _3379_/B vssd1 vssd1 vccd1 vccd1 _3267_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5245_/CLK _5005_/D vssd1 vssd1 vccd1 vccd1 _5005_/Q sky130_fd_sc_hd__dfxtp_1
X_3197_ _3197_/A vssd1 vssd1 vccd1 vccd1 _3285_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5529__119 vssd1 vssd1 vccd1 vccd1 _5529__119/HI _5529__119/LO sky130_fd_sc_hd__conb_1
XFILLER_39_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3120_ _3120_/A vssd1 vssd1 vccd1 vccd1 _3120_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3051_ _3051_/A vssd1 vssd1 vccd1 vccd1 _3126_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5462__52 vssd1 vssd1 vccd1 vccd1 _5462__52/HI _5539_/A sky130_fd_sc_hd__conb_1
XFILLER_16_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3953_ _5264_/Q _3915_/X _3697_/A _3947_/X _3952_/X vssd1 vssd1 vccd1 vccd1 _3953_/X
+ sky130_fd_sc_hd__a2111o_1
X_3884_ hold10/A _3170_/X _3884_/S vssd1 vssd1 vccd1 vccd1 _3885_/A sky130_fd_sc_hd__mux2_1
X_2904_ _2906_/A _2906_/B _2906_/C _2904_/D vssd1 vssd1 vccd1 vccd1 _4964_/A sky130_fd_sc_hd__nor4_4
X_2835_ _2833_/X _5026_/Q _2834_/X vssd1 vssd1 vccd1 vccd1 _2835_/Y sky130_fd_sc_hd__a21oi_1
X_5623_ _5623_/A _2659_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[19] sky130_fd_sc_hd__ebufn_8
X_5554_ _5554_/A _2576_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[20] sky130_fd_sc_hd__ebufn_8
X_2766_ _2766_/A _2766_/B vssd1 vssd1 vccd1 vccd1 _2767_/A sky130_fd_sc_hd__and2_1
X_2697_ _2698_/A vssd1 vssd1 vccd1 vccd1 _2697_/Y sky130_fd_sc_hd__clkinv_4
X_4505_ _5272_/Q _5273_/Q _5271_/Q vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__or3b_1
X_4436_ _4436_/A _4436_/B _4435_/X vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__or3b_1
X_4367_ _4381_/A _4367_/B vssd1 vssd1 vccd1 vccd1 _4367_/X sky130_fd_sc_hd__or2_1
X_3318_ _3318_/A _3318_/B vssd1 vssd1 vccd1 vccd1 _3319_/C sky130_fd_sc_hd__xor2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _4298_/A vssd1 vssd1 vccd1 vccd1 _5215_/D sky130_fd_sc_hd__clkbuf_1
X_3249_ _3247_/B _3247_/C _4953_/B vssd1 vssd1 vccd1 vccd1 _3249_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2620_ _2622_/A vssd1 vssd1 vccd1 vccd1 _2620_/Y sky130_fd_sc_hd__inv_2
X_2551_ _2734_/A _2554_/A _2550_/Y vssd1 vssd1 vccd1 vccd1 _5115_/D sky130_fd_sc_hd__a21oi_1
X_5270_ _5322_/CLK _5270_/D vssd1 vssd1 vccd1 vccd1 _5270_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4221_ _4258_/S vssd1 vssd1 vccd1 vccd1 _4234_/S sky130_fd_sc_hd__clkbuf_2
X_4152_ _4152_/A vssd1 vssd1 vccd1 vccd1 _5176_/D sky130_fd_sc_hd__clkbuf_1
X_4083_ _4083_/A _4083_/B vssd1 vssd1 vccd1 vccd1 _5151_/D sky130_fd_sc_hd__nor2_1
X_3103_ _3118_/S _3115_/B vssd1 vssd1 vccd1 vccd1 _3103_/X sky130_fd_sc_hd__or2_1
XFILLER_55_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3034_ _3035_/A _3035_/B vssd1 vssd1 vccd1 vccd1 _3036_/A sky130_fd_sc_hd__or2_2
XFILLER_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4985_ _5446_/CLK _4985_/D vssd1 vssd1 vccd1 vccd1 _5584_/A sky130_fd_sc_hd__dfxtp_4
X_3936_ _5261_/Q _3919_/X _3897_/X _5083_/Q vssd1 vssd1 vccd1 vccd1 _3936_/X sky130_fd_sc_hd__a22o_1
X_4005__12 _4005__12/A vssd1 vssd1 vccd1 vccd1 _5119_/CLK sky130_fd_sc_hd__inv_2
XFILLER_137_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3867_ hold34/A _4832_/B _3873_/S vssd1 vssd1 vccd1 vccd1 _3868_/A sky130_fd_sc_hd__mux2_1
X_5606_ _5606_/A _2638_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[2] sky130_fd_sc_hd__ebufn_8
X_3798_ _3803_/C _3798_/B _3820_/A vssd1 vssd1 vccd1 vccd1 _3799_/A sky130_fd_sc_hd__and3b_1
X_2818_ _5129_/Q _5130_/Q vssd1 vssd1 vccd1 vccd1 _2822_/B sky130_fd_sc_hd__or2_1
X_5537_ _5537_/A _2686_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[3] sky130_fd_sc_hd__ebufn_8
XFILLER_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2749_ _4634_/A vssd1 vssd1 vccd1 vccd1 _4571_/A sky130_fd_sc_hd__buf_2
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5399_ _5403_/Q _5399_/D vssd1 vssd1 vccd1 vccd1 _5399_/Q sky130_fd_sc_hd__dfxtp_1
X_4419_ _4419_/A _4419_/B vssd1 vssd1 vccd1 vccd1 _4419_/X sky130_fd_sc_hd__or2_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5369_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_23_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput19 la1_data_in[0] vssd1 vssd1 vccd1 vccd1 _4508_/A sky130_fd_sc_hd__buf_6
XFILLER_136_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4770_ _4774_/C _4770_/B vssd1 vssd1 vccd1 vccd1 _5363_/D sky130_fd_sc_hd__nor2_1
X_3721_ _3718_/Y _3720_/X _5017_/Q _3711_/X vssd1 vssd1 vccd1 vccd1 _5017_/D sky130_fd_sc_hd__o2bb2a_1
X_3652_ _3652_/A _3652_/B vssd1 vssd1 vccd1 vccd1 _3653_/S sky130_fd_sc_hd__xnor2_1
X_2603_ _2603_/A vssd1 vssd1 vccd1 vccd1 _2603_/Y sky130_fd_sc_hd__inv_2
X_3583_ _3583_/A _3583_/B vssd1 vssd1 vccd1 vccd1 _4995_/D sky130_fd_sc_hd__nor2_1
X_2534_ _5113_/Q vssd1 vssd1 vccd1 vccd1 _2736_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_5322_ _5322_/CLK _5322_/D vssd1 vssd1 vccd1 vccd1 _5322_/Q sky130_fd_sc_hd__dfxtp_1
X_5253_ _5446_/CLK _5253_/D vssd1 vssd1 vccd1 vccd1 _5253_/Q sky130_fd_sc_hd__dfxtp_1
X_5184_ _5444_/CLK _5184_/D vssd1 vssd1 vccd1 vccd1 _5184_/Q sky130_fd_sc_hd__dfxtp_1
X_4204_ _5414_/Q _5365_/Q _4216_/S vssd1 vssd1 vccd1 vccd1 _4204_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4135_ _5346_/Q _5169_/Q _4137_/S vssd1 vssd1 vccd1 vccd1 _4136_/A sky130_fd_sc_hd__mux2_1
X_4066_ _4066_/A vssd1 vssd1 vccd1 vccd1 _5144_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3017_ _2973_/A _5377_/Q _3016_/X _2980_/A vssd1 vssd1 vccd1 vccd1 _3018_/B sky130_fd_sc_hd__o211a_1
XFILLER_52_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4968_ _4965_/A _4965_/B _5601_/A vssd1 vssd1 vccd1 vccd1 _4968_/X sky130_fd_sc_hd__a21o_1
X_4899_ _5385_/D _4884_/X _4898_/X _4882_/X vssd1 vssd1 vccd1 vccd1 _5417_/D sky130_fd_sc_hd__o211a_1
X_3919_ _3919_/A vssd1 vssd1 vccd1 vccd1 _3919_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_137_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4822_ _4822_/A vssd1 vssd1 vccd1 vccd1 _5400_/D sky130_fd_sc_hd__clkbuf_1
X_4753_ _5358_/Q _4751_/A _4746_/X vssd1 vssd1 vccd1 vccd1 _4754_/B sky130_fd_sc_hd__o21ai_1
X_3704_ _5014_/Q _3697_/X _3700_/X hold141/X vssd1 vssd1 vccd1 vccd1 _5014_/D sky130_fd_sc_hd__a22o_1
X_4684_ _4587_/B _4680_/X _4681_/X _3642_/B vssd1 vssd1 vccd1 vccd1 _4685_/B sky130_fd_sc_hd__o22a_1
X_3635_ _3912_/A _3892_/B vssd1 vssd1 vccd1 vccd1 _3699_/A sky130_fd_sc_hd__nor2_2
X_3566_ _3575_/B _3566_/B _3569_/A vssd1 vssd1 vccd1 vccd1 _3567_/A sky130_fd_sc_hd__and3b_1
X_4002__9 _4002__9/A vssd1 vssd1 vccd1 vccd1 _5116_/CLK sky130_fd_sc_hd__inv_2
X_3497_ _5574_/A _4693_/A vssd1 vssd1 vccd1 vccd1 _3498_/A sky130_fd_sc_hd__and2b_1
X_5305_ _5305_/CLK _5305_/D vssd1 vssd1 vccd1 vccd1 _5305_/Q sky130_fd_sc_hd__dfxtp_1
X_5236_ _5436_/CLK _5236_/D vssd1 vssd1 vccd1 vccd1 _5236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5167_ _5351_/CLK _5167_/D vssd1 vssd1 vccd1 vccd1 _5167_/Q sky130_fd_sc_hd__dfxtp_2
X_4118_ _5338_/Q _5161_/Q _4126_/S vssd1 vssd1 vccd1 vccd1 _4119_/A sky130_fd_sc_hd__mux2_1
X_5098_ _5435_/CLK _5098_/D vssd1 vssd1 vccd1 vccd1 _5098_/Q sky130_fd_sc_hd__dfxtp_1
X_4049_ _4049_/A vssd1 vssd1 vccd1 vccd1 _5136_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3420_ _3417_/X _3418_/X _3420_/S vssd1 vssd1 vccd1 vccd1 _3431_/A sky130_fd_sc_hd__mux2_4
X_3351_ _3344_/X _3350_/X _3267_/A vssd1 vssd1 vccd1 vccd1 _3351_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3282_ _3224_/A _3280_/Y _3281_/X _3279_/B vssd1 vssd1 vccd1 vccd1 _3300_/B sky130_fd_sc_hd__o31ai_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _5058_/CLK _5021_/D vssd1 vssd1 vccd1 vccd1 _5021_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4805_ _4805_/A vssd1 vssd1 vccd1 vccd1 _5392_/D sky130_fd_sc_hd__clkbuf_1
X_2997_ _5307_/Q _2974_/A _2952_/Y input42/X _2892_/A vssd1 vssd1 vccd1 vccd1 _2997_/X
+ sky130_fd_sc_hd__a221o_1
X_4736_ _5337_/Q _5109_/Q _4942_/D vssd1 vssd1 vccd1 vccd1 _4737_/A sky130_fd_sc_hd__and3_1
X_4667_ _4667_/A _4667_/B vssd1 vssd1 vccd1 vccd1 _4668_/A sky130_fd_sc_hd__and2_1
X_3618_ _5322_/Q _5321_/Q vssd1 vssd1 vccd1 vccd1 _3893_/B sky130_fd_sc_hd__nand2_1
X_4598_ _3627_/X _4665_/S _4597_/Y vssd1 vssd1 vccd1 vccd1 _4666_/S sky130_fd_sc_hd__a21oi_4
X_3549_ _3682_/B _3682_/C _3549_/C vssd1 vssd1 vccd1 vccd1 _3549_/X sky130_fd_sc_hd__and3_1
XFILLER_57_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5219_ _5245_/CLK _5219_/D vssd1 vssd1 vccd1 vccd1 _5219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2920_ _5243_/Q vssd1 vssd1 vccd1 vccd1 _4791_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2851_ _5132_/Q vssd1 vssd1 vccd1 vccd1 _4042_/A sky130_fd_sc_hd__buf_2
X_5570_ _5570_/A _2595_/Y vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__ebufn_8
X_2782_ _2782_/A _4092_/A vssd1 vssd1 vccd1 vccd1 _2785_/C sky130_fd_sc_hd__xnor2_1
X_4521_ _4532_/A vssd1 vssd1 vccd1 vccd1 _4530_/S sky130_fd_sc_hd__clkbuf_2
X_4452_ _4455_/B _4450_/Y _4451_/Y _4445_/X _3510_/A vssd1 vssd1 vccd1 vccd1 _4453_/B
+ sky130_fd_sc_hd__o32a_1
X_3403_ _3442_/A _3829_/B _3829_/A _3835_/B vssd1 vssd1 vccd1 vccd1 _3403_/X sky130_fd_sc_hd__a211o_1
X_4383_ _4402_/A vssd1 vssd1 vccd1 vccd1 _4383_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3334_ _3334_/A _3563_/C vssd1 vssd1 vccd1 vccd1 _3357_/A sky130_fd_sc_hd__or2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3265_/A _3265_/B vssd1 vssd1 vccd1 vccd1 _3379_/B sky130_fd_sc_hd__xor2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _5245_/CLK _5004_/D vssd1 vssd1 vccd1 vccd1 _5004_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3196_ _3402_/A _3216_/A _3244_/C _5055_/Q vssd1 vssd1 vccd1 vccd1 _3197_/A sky130_fd_sc_hd__a211o_1
XFILLER_54_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4719_ _5332_/Q _4722_/C vssd1 vssd1 vccd1 vccd1 _4720_/B sky130_fd_sc_hd__or2_1
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5512__102 vssd1 vssd1 vccd1 vccd1 _5512__102/HI _5619_/A sky130_fd_sc_hd__conb_1
XFILLER_13_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3050_ _3108_/A vssd1 vssd1 vccd1 vccd1 _3126_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_23_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3952_ _4553_/A _4594_/B _3912_/A _5086_/Q vssd1 vssd1 vccd1 vccd1 _3952_/X sky130_fd_sc_hd__o31a_1
X_3883_ _3883_/A vssd1 vssd1 vccd1 vccd1 _5074_/D sky130_fd_sc_hd__clkbuf_1
X_2903_ _5372_/Q _2903_/B _2903_/C _2902_/X vssd1 vssd1 vccd1 vccd1 _2904_/D sky130_fd_sc_hd__or4b_1
XFILLER_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2834_ _2795_/X _5025_/Q _3480_/B vssd1 vssd1 vccd1 vccd1 _2834_/X sky130_fd_sc_hd__and3b_1
X_5622_ _5623_/A _2658_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[18] sky130_fd_sc_hd__ebufn_8
X_5553_ _5553_/A _2575_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[19] sky130_fd_sc_hd__ebufn_8
X_2765_ _2760_/A _2768_/A _2768_/B _2764_/X vssd1 vssd1 vccd1 vccd1 _2766_/B sky130_fd_sc_hd__a31o_1
X_4504_ _4504_/A _4504_/B vssd1 vssd1 vccd1 vccd1 _4551_/B sky130_fd_sc_hd__and2_1
X_2696_ _2698_/A vssd1 vssd1 vccd1 vccd1 _2696_/Y sky130_fd_sc_hd__inv_2
X_4435_ _3592_/A _4353_/X _4363_/C _3533_/B vssd1 vssd1 vccd1 vccd1 _4435_/X sky130_fd_sc_hd__o211a_1
X_4366_ input6/X _5161_/Q _4380_/S vssd1 vssd1 vccd1 vccd1 _4367_/B sky130_fd_sc_hd__mux2_1
XFILLER_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3317_ _3751_/A _3424_/A _3409_/A vssd1 vssd1 vccd1 vccd1 _3318_/B sky130_fd_sc_hd__mux2_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4296_/X _5215_/Q _4309_/S vssd1 vssd1 vccd1 vccd1 _4298_/A sky130_fd_sc_hd__mux2_1
X_3248_ _5441_/Q vssd1 vssd1 vccd1 vccd1 _4953_/B sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3179_ _3179_/A _3179_/B vssd1 vssd1 vccd1 vccd1 _3180_/B sky130_fd_sc_hd__and2_1
XFILLER_39_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5508__98 vssd1 vssd1 vccd1 vccd1 _5508__98/HI _5611_/A sky130_fd_sc_hd__conb_1
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2550_ _2734_/A _2554_/A _2530_/B vssd1 vssd1 vccd1 vccd1 _2550_/Y sky130_fd_sc_hd__o21ai_1
X_4220_ _4434_/A _4355_/C _4220_/C vssd1 vssd1 vccd1 vccd1 _4258_/S sky130_fd_sc_hd__and3_2
X_4151_ _5353_/Q _5176_/Q _4180_/S vssd1 vssd1 vccd1 vccd1 _4152_/A sky130_fd_sc_hd__mux2_1
X_4082_ _4084_/B _4092_/B _4081_/X vssd1 vssd1 vccd1 vccd1 _4083_/B sky130_fd_sc_hd__o21ai_1
X_3102_ _3115_/A _3102_/B _3102_/C vssd1 vssd1 vccd1 vccd1 _3102_/X sky130_fd_sc_hd__and3_1
X_3033_ _3033_/A _3033_/B vssd1 vssd1 vccd1 vccd1 _3035_/B sky130_fd_sc_hd__xnor2_2
XFILLER_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4984_ _5446_/CLK _4984_/D vssd1 vssd1 vccd1 vccd1 _5583_/A sky130_fd_sc_hd__dfxtp_4
X_3935_ _5086_/Q _3932_/X _3934_/X vssd1 vssd1 vccd1 vccd1 _5086_/D sky130_fd_sc_hd__o21a_1
X_3866_ _3866_/A vssd1 vssd1 vccd1 vccd1 _5066_/D sky130_fd_sc_hd__clkbuf_1
X_5605_ _5605_/A _2637_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[1] sky130_fd_sc_hd__ebufn_8
X_2817_ _2812_/Y _2815_/Y _2817_/S vssd1 vssd1 vccd1 vccd1 _2817_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3797_ _5044_/Q _3797_/B vssd1 vssd1 vccd1 vccd1 _3798_/B sky130_fd_sc_hd__or2_1
X_5536_ _5536_/A _2683_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[2] sky130_fd_sc_hd__ebufn_8
X_2748_ _4827_/A vssd1 vssd1 vccd1 vccd1 _4634_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2679_ _2683_/A vssd1 vssd1 vccd1 vccd1 _2679_/Y sky130_fd_sc_hd__inv_2
X_4418_ _5205_/Q _5175_/Q _4418_/S vssd1 vssd1 vccd1 vccd1 _4419_/B sky130_fd_sc_hd__mux2_1
X_5398_ _5403_/Q _5398_/D vssd1 vssd1 vccd1 vccd1 _5398_/Q sky130_fd_sc_hd__dfxtp_1
X_4349_ _4349_/A vssd1 vssd1 vccd1 vccd1 _5226_/D sky130_fd_sc_hd__clkbuf_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_136_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3720_ _4038_/A _3720_/B _3729_/B _3736_/A vssd1 vssd1 vccd1 vccd1 _3720_/X sky130_fd_sc_hd__and4b_1
XFILLER_20_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3651_ _5237_/Q _3651_/B vssd1 vssd1 vccd1 vccd1 _3652_/B sky130_fd_sc_hd__nor2_1
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2602_ _2603_/A vssd1 vssd1 vccd1 vccd1 _2602_/Y sky130_fd_sc_hd__inv_2
X_3582_ _4995_/Q _3581_/B _3569_/X vssd1 vssd1 vccd1 vccd1 _3583_/B sky130_fd_sc_hd__o21ai_1
X_2533_ _5115_/Q vssd1 vssd1 vccd1 vccd1 _2734_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5321_ _5322_/CLK _5321_/D vssd1 vssd1 vccd1 vccd1 _5321_/Q sky130_fd_sc_hd__dfxtp_1
X_5499__89 vssd1 vssd1 vccd1 vccd1 _5499__89/HI _5598_/A sky130_fd_sc_hd__conb_1
X_5252_ _5446_/CLK _5252_/D vssd1 vssd1 vccd1 vccd1 _5252_/Q sky130_fd_sc_hd__dfxtp_1
X_5183_ _5444_/CLK _5183_/D vssd1 vssd1 vccd1 vccd1 _5183_/Q sky130_fd_sc_hd__dfxtp_1
X_4203_ _4203_/A vssd1 vssd1 vccd1 vccd1 _4216_/S sky130_fd_sc_hd__clkbuf_2
X_4134_ _4134_/A vssd1 vssd1 vccd1 vccd1 _5168_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4065_ _5381_/Q hold64/A _4065_/S vssd1 vssd1 vccd1 vccd1 _4066_/A sky130_fd_sc_hd__mux2_1
X_3016_ _5308_/Q _3075_/B _2952_/Y input43/X _2975_/A vssd1 vssd1 vccd1 vccd1 _3016_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4967_ _2918_/X _4965_/Y _4966_/X _4902_/X vssd1 vssd1 vccd1 vccd1 _5447_/D sky130_fd_sc_hd__o211a_1
X_4898_ _4900_/B _4897_/X _4884_/A vssd1 vssd1 vccd1 vccd1 _4898_/X sky130_fd_sc_hd__a21bo_1
XFILLER_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3918_ _5081_/Q _3909_/X _3917_/X vssd1 vssd1 vccd1 vccd1 _5081_/D sky130_fd_sc_hd__o21a_1
XFILLER_20_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3849_ _3851_/B _3854_/A _3849_/C vssd1 vssd1 vccd1 vccd1 _3850_/A sky130_fd_sc_hd__and3b_1
XFILLER_20_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4821_ _3170_/X _5400_/Q _4823_/S vssd1 vssd1 vccd1 vccd1 _4822_/A sky130_fd_sc_hd__mux2_1
XFILLER_34_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4752_ _5358_/Q _5357_/Q _4752_/C vssd1 vssd1 vccd1 vccd1 _4758_/C sky130_fd_sc_hd__and3_1
XFILLER_14_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3703_ _5013_/Q _3697_/X _3700_/X _5275_/Q vssd1 vssd1 vccd1 vccd1 _5013_/D sky130_fd_sc_hd__a22o_1
X_4683_ _4328_/B _4680_/X _4681_/X _4682_/X _4350_/X vssd1 vssd1 vccd1 vccd1 _5321_/D
+ sky130_fd_sc_hd__o221a_1
X_3634_ _3626_/Y _3632_/X _3633_/X vssd1 vssd1 vccd1 vccd1 _5000_/D sky130_fd_sc_hd__a21oi_1
X_3565_ _4073_/D _3377_/A _3563_/B _3563_/A vssd1 vssd1 vccd1 vccd1 _3566_/B sky130_fd_sc_hd__a31o_1
X_3496_ _4587_/C vssd1 vssd1 vccd1 vccd1 _4693_/A sky130_fd_sc_hd__clkbuf_2
X_5304_ _5435_/CLK _5304_/D vssd1 vssd1 vccd1 vccd1 _5304_/Q sky130_fd_sc_hd__dfxtp_1
X_5235_ _5436_/CLK _5235_/D vssd1 vssd1 vccd1 vccd1 _5235_/Q sky130_fd_sc_hd__dfxtp_1
X_5166_ _5351_/CLK _5166_/D vssd1 vssd1 vccd1 vccd1 _5166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4117_ _4261_/S vssd1 vssd1 vccd1 vccd1 _4126_/S sky130_fd_sc_hd__clkbuf_2
X_5097_ _5435_/CLK _5097_/D vssd1 vssd1 vccd1 vccd1 _5097_/Q sky130_fd_sc_hd__dfxtp_1
X_4048_ _2902_/X hold58/A _4054_/S vssd1 vssd1 vccd1 vccd1 _4049_/A sky130_fd_sc_hd__mux2_1
XFILLER_56_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_16_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3350_ _3348_/X _3338_/A _3350_/S vssd1 vssd1 vccd1 vccd1 _3350_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3280_/A _3280_/B _3279_/Y vssd1 vssd1 vccd1 vccd1 _3281_/X sky130_fd_sc_hd__o21ba_1
X_5020_ _5058_/CLK _5020_/D vssd1 vssd1 vccd1 vccd1 _5020_/Q sky130_fd_sc_hd__dfxtp_1
X_5469__59 vssd1 vssd1 vccd1 vccd1 _5469__59/HI _5546_/A sky130_fd_sc_hd__conb_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4804_ _4832_/B _5392_/Q _4812_/S vssd1 vssd1 vccd1 vccd1 _4805_/A sky130_fd_sc_hd__mux2_1
X_2996_ _5238_/Q _2996_/B vssd1 vssd1 vccd1 vccd1 _3002_/A sky130_fd_sc_hd__xnor2_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4735_ _5336_/Q _4115_/B _5337_/Q vssd1 vssd1 vccd1 vccd1 _4738_/B sky130_fd_sc_hd__a21oi_1
X_4666_ _5318_/Q _4665_/X _4666_/S vssd1 vssd1 vccd1 vccd1 _4667_/B sky130_fd_sc_hd__mux2_1
X_3617_ _3617_/A vssd1 vssd1 vccd1 vccd1 _3912_/A sky130_fd_sc_hd__clkbuf_2
X_4597_ _3892_/A _3627_/X _4506_/Y _4587_/C vssd1 vssd1 vccd1 vccd1 _4597_/Y sky130_fd_sc_hd__o211ai_2
X_3548_ _5176_/Q _3541_/X _3547_/X _3535_/X vssd1 vssd1 vccd1 vccd1 _3549_/C sky130_fd_sc_hd__a22o_1
X_3479_ _3465_/Y _3475_/X _3478_/X vssd1 vssd1 vccd1 vccd1 _3479_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5218_ _5351_/CLK _5218_/D vssd1 vssd1 vccd1 vccd1 _5218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5149_ _5439_/CLK _5149_/D vssd1 vssd1 vccd1 vccd1 _5149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5483__73 vssd1 vssd1 vccd1 vccd1 _5483__73/HI _5560_/A sky130_fd_sc_hd__conb_1
XFILLER_13_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2850_ _4022_/A vssd1 vssd1 vccd1 vccd1 _3489_/A sky130_fd_sc_hd__clkbuf_2
X_2781_ _5154_/Q _2781_/B vssd1 vssd1 vccd1 vccd1 _4092_/A sky130_fd_sc_hd__and2_1
XFILLER_31_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4520_ _4520_/A vssd1 vssd1 vccd1 vccd1 _5274_/D sky130_fd_sc_hd__clkbuf_1
X_4451_ _4449_/B _4357_/A _5251_/Q vssd1 vssd1 vccd1 vccd1 _4451_/Y sky130_fd_sc_hd__a21oi_1
X_3402_ _3402_/A vssd1 vssd1 vccd1 vccd1 _3835_/B sky130_fd_sc_hd__clkbuf_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4382_ _5232_/Q _4362_/X _4381_/X _4378_/X vssd1 vssd1 vccd1 vccd1 _5232_/D sky130_fd_sc_hd__o211a_1
X_3333_ _4073_/D _4987_/Q vssd1 vssd1 vccd1 vccd1 _3563_/C sky130_fd_sc_hd__and2_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _3264_/A _3225_/X vssd1 vssd1 vccd1 vccd1 _3265_/A sky130_fd_sc_hd__or2b_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5403_/Q _5003_/D vssd1 vssd1 vccd1 vccd1 _5003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3195_ _5060_/Q _5059_/Q _5058_/Q _5057_/Q _5061_/Q vssd1 vssd1 vccd1 vccd1 _3244_/C
+ sky130_fd_sc_hd__a41o_1
XFILLER_38_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2979_ _5454_/Q _4975_/B _2977_/X _2978_/X vssd1 vssd1 vccd1 vccd1 _2979_/X sky130_fd_sc_hd__o211a_1
X_4718_ _5332_/Q _4722_/C vssd1 vssd1 vccd1 vccd1 _4725_/C sky130_fd_sc_hd__and2_1
X_4649_ _5296_/Q _5266_/Q _4661_/S vssd1 vssd1 vccd1 vccd1 _4649_/X sky130_fd_sc_hd__mux2_1
XFILLER_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5431_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_55_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _4587_/A vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2902_ _5373_/Q vssd1 vssd1 vccd1 vccd1 _2902_/X sky130_fd_sc_hd__clkbuf_4
X_3882_ hold19/A _4834_/C _3884_/S vssd1 vssd1 vccd1 vccd1 _3883_/A sky130_fd_sc_hd__mux2_1
XFILLER_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2833_ _2833_/A vssd1 vssd1 vccd1 vccd1 _2833_/X sky130_fd_sc_hd__clkbuf_2
X_5621_ _5623_/A _2657_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[17] sky130_fd_sc_hd__ebufn_8
X_5552_ _5552_/A _2574_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[18] sky130_fd_sc_hd__ebufn_8
X_2764_ _2739_/Y _3754_/A vssd1 vssd1 vccd1 vccd1 _2764_/X sky130_fd_sc_hd__and2b_1
XFILLER_8_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4503_ _5254_/Q _4503_/B vssd1 vssd1 vccd1 vccd1 _4508_/B sky130_fd_sc_hd__nand2_1
X_2695_ _2695_/A vssd1 vssd1 vccd1 vccd1 _2695_/Y sky130_fd_sc_hd__inv_2
X_4434_ _4434_/A _4434_/B _4434_/C vssd1 vssd1 vccd1 vccd1 _4436_/B sky130_fd_sc_hd__and3_1
X_4365_ _4421_/S vssd1 vssd1 vccd1 vccd1 _4380_/S sky130_fd_sc_hd__clkbuf_2
X_3316_ _5061_/Q _3424_/A vssd1 vssd1 vccd1 vccd1 _3751_/A sky130_fd_sc_hd__nor2_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _5211_/Q _4275_/X _4295_/X vssd1 vssd1 vccd1 vccd1 _4296_/X sky130_fd_sc_hd__a21o_1
X_3247_ _5441_/Q _3247_/B _3247_/C vssd1 vssd1 vccd1 vccd1 _3250_/A sky130_fd_sc_hd__and3_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _3179_/A _3179_/B vssd1 vssd1 vccd1 vccd1 _3646_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4150_ _4200_/A vssd1 vssd1 vccd1 vccd1 _4180_/S sky130_fd_sc_hd__clkbuf_2
X_3101_ _3115_/A _3102_/B _3102_/C vssd1 vssd1 vccd1 vccd1 _3101_/Y sky130_fd_sc_hd__a21oi_1
X_4081_ _4350_/A vssd1 vssd1 vccd1 vccd1 _4081_/X sky130_fd_sc_hd__clkbuf_2
X_5519__109 vssd1 vssd1 vccd1 vccd1 _5519__109/HI _5635_/A sky130_fd_sc_hd__conb_1
X_3032_ _2973_/A _5378_/Q _3031_/X _2980_/A vssd1 vssd1 vccd1 vccd1 _3033_/B sky130_fd_sc_hd__o211a_1
XFILLER_36_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4983_ _5454_/Q _4980_/B _4982_/X _4861_/A vssd1 vssd1 vccd1 vccd1 _5454_/D sky130_fd_sc_hd__o211a_1
XFILLER_23_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3934_ _5082_/Q _3904_/C _3933_/X _3911_/X vssd1 vssd1 vccd1 vccd1 _3934_/X sky130_fd_sc_hd__a211o_1
X_3865_ hold25/A _4832_/A _3873_/S vssd1 vssd1 vccd1 vccd1 _3866_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5604_ _5604_/A _2697_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[0] sky130_fd_sc_hd__ebufn_8
X_2816_ _5130_/Q _2816_/B vssd1 vssd1 vccd1 vccd1 _2817_/S sky130_fd_sc_hd__xnor2_2
X_3796_ _5044_/Q _3797_/B vssd1 vssd1 vccd1 vccd1 _3803_/C sky130_fd_sc_hd__and2_1
XFILLER_11_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5535_ _5535_/A _2685_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[1] sky130_fd_sc_hd__ebufn_8
X_2747_ _4158_/A vssd1 vssd1 vccd1 vccd1 _4827_/A sky130_fd_sc_hd__buf_4
X_2678_ _2690_/A vssd1 vssd1 vccd1 vccd1 _2683_/A sky130_fd_sc_hd__buf_8
X_4417_ _5241_/Q _4402_/X _4415_/X _4416_/X vssd1 vssd1 vccd1 vccd1 _5241_/D sky130_fd_sc_hd__o211a_1
X_5397_ _5403_/Q _5397_/D vssd1 vssd1 vccd1 vccd1 _5397_/Q sky130_fd_sc_hd__dfxtp_1
X_4348_ _4348_/A _4348_/B vssd1 vssd1 vccd1 vccd1 _4349_/A sky130_fd_sc_hd__or2_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4279_ _4278_/X _5211_/Q _4288_/S vssd1 vssd1 vccd1 vccd1 _4280_/A sky130_fd_sc_hd__mux2_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3650_ _5318_/Q _3076_/X _3645_/Y _3155_/B vssd1 vssd1 vccd1 vccd1 _3651_/B sky130_fd_sc_hd__o2bb2a_1
X_2601_ _2603_/A vssd1 vssd1 vccd1 vccd1 _2601_/Y sky130_fd_sc_hd__inv_2
X_3581_ _4995_/Q _3581_/B vssd1 vssd1 vccd1 vccd1 _3583_/A sky130_fd_sc_hd__and2_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5320_ _5435_/CLK _5320_/D vssd1 vssd1 vccd1 vccd1 _5320_/Q sky130_fd_sc_hd__dfxtp_4
X_2532_ _5118_/Q vssd1 vssd1 vccd1 vccd1 _3705_/A sky130_fd_sc_hd__clkbuf_2
X_5251_ _5446_/CLK _5251_/D vssd1 vssd1 vccd1 vccd1 _5251_/Q sky130_fd_sc_hd__dfxtp_1
X_4202_ _4202_/A vssd1 vssd1 vccd1 vccd1 _5189_/D sky130_fd_sc_hd__clkbuf_1
X_5182_ _5339_/CLK _5182_/D vssd1 vssd1 vccd1 vccd1 _5182_/Q sky130_fd_sc_hd__dfxtp_1
X_4133_ _5345_/Q _5168_/Q _4137_/S vssd1 vssd1 vccd1 vccd1 _4134_/A sky130_fd_sc_hd__mux2_1
X_4064_ _4064_/A vssd1 vssd1 vccd1 vccd1 _5143_/D sky130_fd_sc_hd__clkbuf_1
X_3015_ _3051_/A _3015_/B vssd1 vssd1 vccd1 vccd1 _3020_/A sky130_fd_sc_hd__xnor2_1
XFILLER_36_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4966_ _4965_/A _4965_/B _5600_/A vssd1 vssd1 vccd1 vccd1 _4966_/X sky130_fd_sc_hd__a21o_1
X_4897_ _5417_/Q _4897_/B vssd1 vssd1 vccd1 vccd1 _4897_/X sky130_fd_sc_hd__or2_1
X_3917_ _5281_/Q _3910_/X _3911_/X _3916_/X vssd1 vssd1 vccd1 vccd1 _3917_/X sky130_fd_sc_hd__a211o_1
X_3848_ _3835_/A _3749_/B _3834_/A _3824_/B vssd1 vssd1 vccd1 vccd1 _3849_/C sky130_fd_sc_hd__a31o_1
X_3779_ _3729_/A _3779_/A2 _3764_/S _3230_/Y _3750_/X vssd1 vssd1 vccd1 vccd1 _3779_/X
+ sky130_fd_sc_hd__a32o_1
X_5449_ _5403_/Q _5449_/D vssd1 vssd1 vccd1 vccd1 _5602_/A sky130_fd_sc_hd__dfxtp_4
XFILLER_28_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4820_ _4820_/A vssd1 vssd1 vccd1 vccd1 _5399_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4751_ _4751_/A _4751_/B vssd1 vssd1 vccd1 vccd1 _5357_/D sky130_fd_sc_hd__nor2_1
X_3702_ _5012_/Q _3697_/X _3700_/X _5276_/Q vssd1 vssd1 vccd1 vccd1 _5012_/D sky130_fd_sc_hd__a22o_1
X_4682_ _5301_/Q _3894_/B _4464_/C vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__a21o_1
X_3633_ _3891_/B _3643_/S _5000_/Q vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__o21ba_1
X_3564_ _3578_/C vssd1 vssd1 vccd1 vccd1 _3575_/B sky130_fd_sc_hd__clkbuf_1
X_5303_ _5435_/CLK _5303_/D vssd1 vssd1 vccd1 vccd1 _5303_/Q sky130_fd_sc_hd__dfxtp_1
X_3495_ _5254_/Q vssd1 vssd1 vccd1 vccd1 _4587_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_5234_ _5436_/CLK _5234_/D vssd1 vssd1 vccd1 vccd1 _5234_/Q sky130_fd_sc_hd__dfxtp_1
X_5165_ _5351_/CLK _5165_/D vssd1 vssd1 vccd1 vccd1 _5165_/Q sky130_fd_sc_hd__dfxtp_1
X_4116_ _4200_/A vssd1 vssd1 vccd1 vccd1 _4261_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_56_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5096_ _5305_/CLK _5096_/D vssd1 vssd1 vccd1 vccd1 _5096_/Q sky130_fd_sc_hd__dfxtp_1
X_4047_ _4047_/A vssd1 vssd1 vccd1 vccd1 _5135_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4949_ _4953_/C _4949_/B vssd1 vssd1 vccd1 vccd1 _5440_/D sky130_fd_sc_hd__nor2_1
XFILLER_24_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3280_ _3280_/A _3280_/B _3279_/Y vssd1 vssd1 vccd1 vccd1 _3280_/Y sky130_fd_sc_hd__nor3b_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4803_ _4825_/S vssd1 vssd1 vccd1 vccd1 _4812_/S sky130_fd_sc_hd__clkbuf_2
X_2995_ _3029_/A _5391_/Q vssd1 vssd1 vccd1 vccd1 _2996_/B sky130_fd_sc_hd__and2_1
X_4734_ _4734_/A vssd1 vssd1 vccd1 vccd1 _5336_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4665_ _5300_/Q _5270_/Q _4665_/S vssd1 vssd1 vccd1 vccd1 _4665_/X sky130_fd_sc_hd__mux2_1
X_4596_ input2/X _5255_/Q _4616_/S vssd1 vssd1 vccd1 vccd1 _4596_/X sky130_fd_sc_hd__mux2_1
X_3616_ _5000_/Q _5001_/Q _5002_/Q vssd1 vssd1 vccd1 vccd1 _3617_/A sky130_fd_sc_hd__or3b_1
X_3547_ _5222_/Q _3547_/B vssd1 vssd1 vccd1 vccd1 _3547_/X sky130_fd_sc_hd__or2_1
X_3478_ _2813_/Y _2814_/X _3476_/Y _3477_/X vssd1 vssd1 vccd1 vccd1 _3478_/X sky130_fd_sc_hd__o211a_1
X_5217_ _5369_/CLK _5217_/D vssd1 vssd1 vccd1 vccd1 _5217_/Q sky130_fd_sc_hd__dfxtp_1
X_5148_ _5328_/CLK _5148_/D vssd1 vssd1 vccd1 vccd1 _5148_/Q sky130_fd_sc_hd__dfxtp_1
X_5079_ _5431_/CLK _5079_/D vssd1 vssd1 vccd1 vccd1 _5079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2780_ _2780_/A _2781_/B vssd1 vssd1 vccd1 vccd1 _2785_/B sky130_fd_sc_hd__xnor2_1
XFILLER_8_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4450_ _4450_/A _4450_/B vssd1 vssd1 vccd1 vccd1 _4450_/Y sky130_fd_sc_hd__nand2_1
X_3401_ _5055_/Q vssd1 vssd1 vccd1 vccd1 _3835_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4381_ _4381_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4381_/X sky130_fd_sc_hd__or2_1
X_3332_ _4989_/Q vssd1 vssd1 vccd1 vccd1 _3551_/B sky130_fd_sc_hd__clkbuf_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _3263_/A _3263_/B vssd1 vssd1 vccd1 vccd1 _3393_/A sky130_fd_sc_hd__xnor2_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ _5053_/Q vssd1 vssd1 vccd1 vccd1 _3216_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5323_/CLK _5002_/D vssd1 vssd1 vccd1 vccd1 _5002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2978_ _5603_/A _4964_/A _2953_/C vssd1 vssd1 vccd1 vccd1 _2978_/X sky130_fd_sc_hd__a21o_1
X_4717_ _4717_/A vssd1 vssd1 vccd1 vccd1 _5331_/D sky130_fd_sc_hd__clkbuf_1
X_4648_ _4648_/A vssd1 vssd1 vccd1 vccd1 _5313_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4579_ _5299_/Q _4581_/B vssd1 vssd1 vccd1 vccd1 _4579_/X sky130_fd_sc_hd__or2_1
XFILLER_45_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3950_ _5089_/Q _3932_/X _3949_/X vssd1 vssd1 vccd1 vccd1 _5089_/D sky130_fd_sc_hd__o21a_1
XFILLER_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2901_ _5374_/Q vssd1 vssd1 vccd1 vccd1 _2903_/C sky130_fd_sc_hd__clkbuf_4
X_3881_ _3881_/A vssd1 vssd1 vccd1 vccd1 _5073_/D sky130_fd_sc_hd__clkbuf_1
X_2832_ _3466_/A _3466_/B vssd1 vssd1 vccd1 vccd1 _2832_/X sky130_fd_sc_hd__or2_1
X_5620_ _5623_/A _2656_/Y vssd1 vssd1 vccd1 vccd1 io_oeb[16] sky130_fd_sc_hd__ebufn_8
X_2763_ _4634_/A vssd1 vssd1 vccd1 vccd1 _2766_/A sky130_fd_sc_hd__buf_4
X_5551_ _5551_/A _2572_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[17] sky130_fd_sc_hd__ebufn_8
XFILLER_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4502_ _4502_/A vssd1 vssd1 vccd1 vccd1 _5270_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2694_ _2695_/A vssd1 vssd1 vccd1 vccd1 _2694_/Y sky130_fd_sc_hd__inv_2
X_4433_ _4433_/A vssd1 vssd1 vccd1 vccd1 _4438_/A sky130_fd_sc_hd__inv_2
X_4364_ _4422_/A vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__clkbuf_1
X_3315_ _3388_/A _3388_/B _3412_/B _3314_/X vssd1 vssd1 vccd1 vccd1 _3319_/B sky130_fd_sc_hd__a211o_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4295_ _5165_/Q _4285_/X _4276_/X _5191_/Q vssd1 vssd1 vccd1 vccd1 _4295_/X sky130_fd_sc_hd__a22o_1
X_3246_ _3221_/B _3221_/C _3221_/A vssd1 vssd1 vccd1 vccd1 _3251_/A sky130_fd_sc_hd__a21bo_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _3652_/A _3177_/B vssd1 vssd1 vccd1 vccd1 _3179_/B sky130_fd_sc_hd__xnor2_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3100_ _3115_/B _3100_/B vssd1 vssd1 vccd1 vccd1 _3102_/C sky130_fd_sc_hd__nand2_1
X_4080_ _4080_/A vssd1 vssd1 vccd1 vccd1 _4092_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3031_ _5309_/Q _2974_/A _2952_/Y input44/X _2975_/A vssd1 vssd1 vccd1 vccd1 _3031_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_36_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4982_ _4982_/A _4982_/B vssd1 vssd1 vccd1 vccd1 _4982_/X sky130_fd_sc_hd__or2_1
XFILLER_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3933_ _5260_/Q _3919_/X _3910_/A _5286_/Q vssd1 vssd1 vccd1 vccd1 _3933_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_3_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5132_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3864_ _3888_/S vssd1 vssd1 vccd1 vccd1 _3873_/S sky130_fd_sc_hd__clkbuf_2
X_5603_ _5603_/A _2636_/Y vssd1 vssd1 vccd1 vccd1 io_out[37] sky130_fd_sc_hd__ebufn_8
X_2815_ _4999_/Q _2813_/B _2813_/Y _2814_/X vssd1 vssd1 vccd1 vccd1 _2815_/Y sky130_fd_sc_hd__a22oi_1
X_3795_ _3795_/A vssd1 vssd1 vccd1 vccd1 _5043_/D sky130_fd_sc_hd__clkbuf_1
X_5534_ _5534_/A _2691_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[0] sky130_fd_sc_hd__ebufn_8
X_2746_ _4508_/A vssd1 vssd1 vccd1 vccd1 _4158_/A sky130_fd_sc_hd__inv_2
X_2677_ _2677_/A vssd1 vssd1 vccd1 vccd1 _2677_/Y sky130_fd_sc_hd__inv_2
X_4416_ _4571_/A vssd1 vssd1 vccd1 vccd1 _4416_/X sky130_fd_sc_hd__clkbuf_4
X_5396_ _5403_/Q _5396_/D vssd1 vssd1 vccd1 vccd1 _5396_/Q sky130_fd_sc_hd__dfxtp_1
X_4347_ _5579_/A _4346_/X _4347_/S vssd1 vssd1 vccd1 vccd1 _4348_/B sky130_fd_sc_hd__mux2_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4278_ _5007_/Q _4275_/X _4277_/X vssd1 vssd1 vccd1 vccd1 _4278_/X sky130_fd_sc_hd__a21o_1
X_3229_ _3285_/B _3229_/B _3229_/C vssd1 vssd1 vccd1 vccd1 _3252_/S sky130_fd_sc_hd__and3_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2600_ _2603_/A vssd1 vssd1 vccd1 vccd1 _2600_/Y sky130_fd_sc_hd__inv_2
X_3580_ _3581_/B _3580_/B vssd1 vssd1 vccd1 vccd1 _4994_/D sky130_fd_sc_hd__nor2_1
X_2531_ _2531_/A vssd1 vssd1 vccd1 vccd1 _5119_/D sky130_fd_sc_hd__clkbuf_1
X_5250_ _5446_/CLK _5250_/D vssd1 vssd1 vccd1 vccd1 _5250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4201_ _4199_/X _5189_/Q _4214_/S vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__mux2_1
X_5181_ _5339_/CLK _5181_/D vssd1 vssd1 vccd1 vccd1 _5181_/Q sky130_fd_sc_hd__dfxtp_1
X_4132_ _4132_/A vssd1 vssd1 vccd1 vccd1 _5167_/D sky130_fd_sc_hd__clkbuf_1
X_4063_ _5380_/Q hold85/A _4065_/S vssd1 vssd1 vccd1 vccd1 _4064_/A sky130_fd_sc_hd__mux2_1
X_3014_ _3029_/A _5392_/Q vssd1 vssd1 vccd1 vccd1 _3015_/B sky130_fd_sc_hd__and2_1
XFILLER_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4965_ _4965_/A _4965_/B vssd1 vssd1 vccd1 vccd1 _4965_/Y sky130_fd_sc_hd__nand2_1
X_3916_ _5255_/Q _3915_/X _3904_/C _5011_/Q vssd1 vssd1 vccd1 vccd1 _3916_/X sky130_fd_sc_hd__a22o_1
X_4896_ _5417_/Q _4897_/B vssd1 vssd1 vccd1 vccd1 _4900_/B sky130_fd_sc_hd__nand2_1
XFILLER_22_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3847_ _3847_/A _3847_/B _3847_/C vssd1 vssd1 vccd1 vccd1 _3851_/B sky130_fd_sc_hd__and3_1
XFILLER_137_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ _3778_/A vssd1 vssd1 vccd1 vccd1 _5031_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2729_ _3705_/C _3705_/D _2729_/C vssd1 vssd1 vccd1 vccd1 _3752_/A sky130_fd_sc_hd__nor3_1
X_5448_ _5403_/Q _5448_/D vssd1 vssd1 vccd1 vccd1 _5601_/A sky130_fd_sc_hd__dfxtp_4
X_5379_ _5403_/Q _5379_/D vssd1 vssd1 vccd1 vccd1 _5379_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4750_ _5357_/Q _4752_/C _4746_/X vssd1 vssd1 vccd1 vccd1 _4751_/B sky130_fd_sc_hd__o21ai_1
XFILLER_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3701_ _5011_/Q _3697_/X _3700_/X _5277_/Q vssd1 vssd1 vccd1 vccd1 _5011_/D sky130_fd_sc_hd__a22o_1
X_4681_ _4681_/A _4680_/X vssd1 vssd1 vccd1 vccd1 _4681_/X sky130_fd_sc_hd__or2b_1
X_3632_ _3912_/B _3627_/X _3892_/B _3631_/Y _5000_/Q vssd1 vssd1 vccd1 vccd1 _3632_/X
+ sky130_fd_sc_hd__a32o_1
X_3563_ _3563_/A _3563_/B _3563_/C vssd1 vssd1 vccd1 vccd1 _3578_/C sky130_fd_sc_hd__and3_1
X_5302_ _5328_/CLK _5302_/D vssd1 vssd1 vccd1 vccd1 _5302_/Q sky130_fd_sc_hd__dfxtp_2
X_3494_ _3494_/A vssd1 vssd1 vccd1 vccd1 _5581_/A sky130_fd_sc_hd__clkbuf_1
X_5233_ _5445_/CLK _5233_/D vssd1 vssd1 vccd1 vccd1 _5233_/Q sky130_fd_sc_hd__dfxtp_1
X_5164_ _5339_/CLK _5164_/D vssd1 vssd1 vccd1 vccd1 _5164_/Q sky130_fd_sc_hd__dfxtp_1
X_4115_ _4115_/A _4115_/B _4436_/A vssd1 vssd1 vccd1 vccd1 _4200_/A sky130_fd_sc_hd__or3_4
XFILLER_29_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5095_ _5305_/CLK _5095_/D vssd1 vssd1 vccd1 vccd1 _5095_/Q sky130_fd_sc_hd__dfxtp_1
X_4046_ _2977_/A hold55/A _4054_/S vssd1 vssd1 vccd1 vccd1 _4047_/A sky130_fd_sc_hd__mux2_1
X_3997__5 _3999__7/A vssd1 vssd1 vccd1 vccd1 _5112_/CLK sky130_fd_sc_hd__inv_2
XFILLER_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4948_ _5440_/Q _4947_/B _2766_/A vssd1 vssd1 vccd1 vccd1 _4949_/B sky130_fd_sc_hd__o21ai_1
XFILLER_33_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4879_ _5413_/Q _4880_/B vssd1 vssd1 vccd1 vccd1 _4888_/C sky130_fd_sc_hd__and2_1
XFILLER_4_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2994_ _2994_/A vssd1 vssd1 vccd1 vccd1 _3041_/A sky130_fd_sc_hd__clkbuf_2
X_4802_ _4802_/A vssd1 vssd1 vccd1 vccd1 _5391_/D sky130_fd_sc_hd__clkbuf_1
X_4733_ _4789_/B _4942_/D _4733_/C vssd1 vssd1 vccd1 vccd1 _4734_/A sky130_fd_sc_hd__and3_1
XFILLER_30_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4664_ _4664_/A vssd1 vssd1 vccd1 vccd1 _5317_/D sky130_fd_sc_hd__clkbuf_1
X_4595_ _4665_/S vssd1 vssd1 vccd1 vccd1 _4616_/S sky130_fd_sc_hd__buf_2
X_3615_ _4594_/A _4587_/B _4594_/B vssd1 vssd1 vccd1 vccd1 _3946_/A sky130_fd_sc_hd__a21o_1
X_3546_ _5584_/A _3677_/B _3545_/X _2761_/X vssd1 vssd1 vccd1 vccd1 _4985_/D sky130_fd_sc_hd__a211o_1
X_3477_ _2846_/A _4999_/Q _3466_/A vssd1 vssd1 vccd1 vccd1 _3477_/X sky130_fd_sc_hd__a21o_1
X_5216_ _5339_/CLK _5216_/D vssd1 vssd1 vccd1 vccd1 _5216_/Q sky130_fd_sc_hd__dfxtp_1
X_5147_ _5313_/CLK _5147_/D vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5078_ _5431_/CLK _5078_/D vssd1 vssd1 vccd1 vccd1 _5078_/Q sky130_fd_sc_hd__dfxtp_1
X_4029_ _3489_/A _2813_/B _4022_/B _4028_/X _4025_/Y vssd1 vssd1 vccd1 vccd1 _5128_/D
+ sky130_fd_sc_hd__a311o_1
XFILLER_13_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5474__64 vssd1 vssd1 vccd1 vccd1 _5474__64/HI _5551_/A sky130_fd_sc_hd__conb_1
XFILLER_16_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3400_ _3424_/C vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4380_ _5195_/Q _5165_/Q _4380_/S vssd1 vssd1 vccd1 vccd1 _4381_/B sky130_fd_sc_hd__mux2_1
X_3331_ _3344_/A _3380_/A _3341_/B vssd1 vssd1 vccd1 vccd1 _3390_/A sky130_fd_sc_hd__or3_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3309_/A _3309_/B vssd1 vssd1 vccd1 vccd1 _3263_/B sky130_fd_sc_hd__xnor2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _5054_/Q vssd1 vssd1 vccd1 vccd1 _3402_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5323_/CLK _5001_/D vssd1 vssd1 vccd1 vccd1 _5001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2977_ _2977_/A _2977_/B _2977_/C vssd1 vssd1 vccd1 vccd1 _2977_/X sky130_fd_sc_hd__or3_1
X_4716_ _4722_/C _4716_/B _4720_/C vssd1 vssd1 vccd1 vccd1 _4717_/A sky130_fd_sc_hd__and3b_1
X_4647_ _4655_/A _4647_/B vssd1 vssd1 vccd1 vccd1 _4648_/A sky130_fd_sc_hd__and2_1
X_4578_ _5294_/Q _4566_/X _4577_/X _4571_/X vssd1 vssd1 vccd1 vccd1 _5298_/D sky130_fd_sc_hd__o211a_1
X_3529_ _3529_/A _3658_/B vssd1 vssd1 vccd1 vccd1 _3547_/B sky130_fd_sc_hd__and2_1
XFILLER_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_0_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5351_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__clkbuf_2
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2900_ _5375_/Q vssd1 vssd1 vccd1 vccd1 _2903_/B sky130_fd_sc_hd__clkbuf_4
X_3880_ hold28/A _4833_/C _3884_/S vssd1 vssd1 vccd1 vccd1 _3881_/A sky130_fd_sc_hd__mux2_1
X_2831_ _2795_/X _5024_/Q _3480_/B _2830_/X _5023_/Q vssd1 vssd1 vccd1 vccd1 _3466_/B
+ sky130_fd_sc_hd__a32o_1
X_5550_ _5550_/A _2571_/Y vssd1 vssd1 vccd1 vccd1 la1_data_out[16] sky130_fd_sc_hd__ebufn_8
X_2762_ _2759_/X _2760_/Y _2761_/X vssd1 vssd1 vccd1 vccd1 _5040_/D sky130_fd_sc_hd__a21oi_1
X_4501_ _5270_/Q _5108_/Q _4519_/S vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__mux2_1
X_2693_ _2695_/A vssd1 vssd1 vccd1 vccd1 _2693_/Y sky130_fd_sc_hd__inv_2
XANTENNA_0 _3420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4432_ _4432_/A vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4363_ _4739_/A _4363_/B _4363_/C vssd1 vssd1 vccd1 vccd1 _4422_/A sky130_fd_sc_hd__nand3_2
X_3314_ _3314_/A _3314_/B vssd1 vssd1 vccd1 vccd1 _3314_/X sky130_fd_sc_hd__and2_1
X_4294_ _4294_/A vssd1 vssd1 vccd1 vccd1 _5214_/D sky130_fd_sc_hd__clkbuf_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3247_/B _3247_/C vssd1 vssd1 vccd1 vccd1 _3245_/X sky130_fd_sc_hd__and2_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _3176_/A _3176_/B vssd1 vssd1 vccd1 vccd1 _3177_/B sky130_fd_sc_hd__and2_1
XFILLER_54_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_136_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3030_ _3051_/A _3030_/B vssd1 vssd1 vccd1 vccd1 _3035_/A sky130_fd_sc_hd__xnor2_1
XFILLER_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4981_ input17/X _4982_/B _4980_/X _4861_/A vssd1 vssd1 vccd1 vccd1 _5453_/D sky130_fd_sc_hd__o211a_1
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3932_ _3956_/S vssd1 vssd1 vccd1 vccd1 _3932_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3863_ _3863_/A vssd1 vssd1 vccd1 vccd1 _5065_/D sky130_fd_sc_hd__clkbuf_1
X_5602_ _5602_/A _2634_/Y vssd1 vssd1 vccd1 vccd1 io_out[36] sky130_fd_sc_hd__ebufn_8
X_2814_ _5035_/Q _4998_/Q _2869_/A vssd1 vssd1 vccd1 vccd1 _2814_/X sky130_fd_sc_hd__mux2_1
X_3794_ _3797_/B _3794_/B _3820_/A vssd1 vssd1 vccd1 vccd1 _3795_/A sky130_fd_sc_hd__and3b_1
X_2745_ _3750_/A _2759_/A _2739_/Y _3729_/A _2744_/X vssd1 vssd1 vccd1 vccd1 _2745_/X
+ sky130_fd_sc_hd__a221o_1
X_2676_ _2677_/A vssd1 vssd1 vccd1 vccd1 _2676_/Y sky130_fd_sc_hd__inv_2
X_5395_ _5403_/Q _5395_/D vssd1 vssd1 vccd1 vccd1 _5395_/Q sky130_fd_sc_hd__dfxtp_1
X_4415_ _4419_/A _4415_/B vssd1 vssd1 vccd1 vccd1 _4415_/X sky130_fd_sc_hd__or2_1
X_4346_ _5270_/Q _3919_/A _3943_/A _5092_/Q _3947_/A vssd1 vssd1 vccd1 vccd1 _4346_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4277_ _5161_/Q _3541_/X _4276_/X _5187_/Q vssd1 vssd1 vccd1 vccd1 _4277_/X sky130_fd_sc_hd__a22o_1
X_3228_ _3402_/A _3216_/A _3823_/D _3284_/A _3205_/Y vssd1 vssd1 vccd1 vccd1 _3229_/C
+ sky130_fd_sc_hd__a41oi_2
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3159_ _3074_/X _2889_/B _3076_/X _5316_/Q vssd1 vssd1 vccd1 vccd1 _3160_/B sky130_fd_sc_hd__a22o_1
XFILLER_27_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2530_ _2527_/B _2530_/B vssd1 vssd1 vccd1 vccd1 _2531_/A sky130_fd_sc_hd__and2b_1
X_5525__115 vssd1 vssd1 vccd1 vccd1 _5525__115/HI _5641_/A sky130_fd_sc_hd__conb_1
X_4200_ _4200_/A vssd1 vssd1 vccd1 vccd1 _4214_/S sky130_fd_sc_hd__clkbuf_2
X_5180_ _5444_/CLK _5180_/D vssd1 vssd1 vccd1 vccd1 _5180_/Q sky130_fd_sc_hd__dfxtp_1
X_4131_ _5344_/Q _5167_/Q _4137_/S vssd1 vssd1 vccd1 vccd1 _4132_/A sky130_fd_sc_hd__mux2_1
X_4062_ _4062_/A vssd1 vssd1 vccd1 vccd1 _5142_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_56_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3013_ _3041_/A _3013_/B _3013_/C vssd1 vssd1 vccd1 vccd1 _3024_/A sky130_fd_sc_hd__and3_1
XFILLER_36_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4964_ _4964_/A vssd1 vssd1 vccd1 vccd1 _4965_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3915_ _3915_/A vssd1 vssd1 vccd1 vccd1 _3915_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4895_ _5384_/D _4884_/X _4894_/Y _4882_/X vssd1 vssd1 vccd1 vccd1 _5416_/D sky130_fd_sc_hd__o211a_1
XFILLER_137_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3846_ _3824_/C _3841_/X _3845_/Y vssd1 vssd1 vccd1 vccd1 _5058_/D sky130_fd_sc_hd__a21oi_1
X_3777_ _3776_/X _5031_/Q _3780_/S vssd1 vssd1 vccd1 vccd1 _3778_/A sky130_fd_sc_hd__mux2_1
X_2728_ _2760_/C _2768_/B _5150_/Q _5038_/Q vssd1 vssd1 vccd1 vccd1 _2728_/X sky130_fd_sc_hd__and4bb_1
X_5447_ _5403_/Q _5447_/D vssd1 vssd1 vccd1 vccd1 _5600_/A sky130_fd_sc_hd__dfxtp_4
X_2659_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2659_/Y sky130_fd_sc_hd__inv_2
X_5378_ _5403_/Q _5378_/D vssd1 vssd1 vccd1 vccd1 _5378_/Q sky130_fd_sc_hd__dfxtp_4
X_4329_ _5089_/Q _3946_/B _4681_/A _4553_/A vssd1 vssd1 vccd1 vccd1 _4329_/X sky130_fd_sc_hd__o211a_1
XFILLER_47_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_136_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_136_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3700_ _4611_/A _3910_/A _4347_/S vssd1 vssd1 vccd1 vccd1 _3700_/X sky130_fd_sc_hd__and3_2
X_4680_ _4678_/X _4680_/B _4680_/C _4680_/D vssd1 vssd1 vccd1 vccd1 _4680_/X sky130_fd_sc_hd__and4b_1
X_3631_ _3642_/A _3891_/B vssd1 vssd1 vccd1 vccd1 _3631_/Y sky130_fd_sc_hd__nor2_1
X_3562_ _3563_/B _3563_/C _3561_/Y vssd1 vssd1 vccd1 vccd1 _4989_/D sky130_fd_sc_hd__a21oi_1
X_5301_ _5323_/CLK _5301_/D vssd1 vssd1 vccd1 vccd1 _5301_/Q sky130_fd_sc_hd__dfxtp_1
X_3493_ _5580_/A _4739_/A vssd1 vssd1 vccd1 vccd1 _3494_/A sky130_fd_sc_hd__and2b_2
X_5232_ _5445_/CLK _5232_/D vssd1 vssd1 vccd1 vccd1 _5232_/Q sky130_fd_sc_hd__dfxtp_1
X_5163_ _5339_/CLK _5163_/D vssd1 vssd1 vccd1 vccd1 _5163_/Q sky130_fd_sc_hd__dfxtp_1
X_4114_ _4115_/B _4113_/X _4355_/C vssd1 vssd1 vccd1 vccd1 _4436_/A sky130_fd_sc_hd__o21ai_1
XFILLER_29_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5094_ _5305_/CLK _5094_/D vssd1 vssd1 vccd1 vccd1 _5094_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4045_ _4071_/S vssd1 vssd1 vccd1 vccd1 _4054_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4947_ _5440_/Q _4947_/B vssd1 vssd1 vccd1 vccd1 _4953_/C sky130_fd_sc_hd__and2_1
X_4878_ _5380_/D _4863_/X _4877_/Y _4861_/X vssd1 vssd1 vccd1 vccd1 _5412_/D sky130_fd_sc_hd__o211a_1
XFILLER_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_137_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3829_ _3829_/A _3829_/B _3829_/C vssd1 vssd1 vccd1 vccd1 _3835_/C sky130_fd_sc_hd__and3_1
XFILLER_28_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_137_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4801_ _4832_/A _5391_/Q _4801_/S vssd1 vssd1 vccd1 vccd1 _4802_/A sky130_fd_sc_hd__mux2_1
X_2993_ _3023_/A vssd1 vssd1 vccd1 vccd1 _3134_/A sky130_fd_sc_hd__buf_6
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4732_ _4789_/A _5227_/Q _4945_/C _4731_/Y _5336_/Q vssd1 vssd1 vccd1 vccd1 _4733_/C
+ sky130_fd_sc_hd__a41o_1
X_4663_ _4667_/A _4663_/B vssd1 vssd1 vccd1 vccd1 _4664_/A sky130_fd_sc_hd__and2_1
X_3614_ _4504_/B vssd1 vssd1 vccd1 vccd1 _4594_/B sky130_fd_sc_hd__clkbuf_2
X_4594_ _4594_/A _4594_/B vssd1 vssd1 vccd1 vccd1 _4665_/S sky130_fd_sc_hd__nand2_4
X_3545_ _3682_/B _3682_/C _3545_/C vssd1 vssd1 vccd1 vccd1 _3545_/X sky130_fd_sc_hd__and3_1
X_3476_ _3476_/A _3476_/B vssd1 vssd1 vccd1 vccd1 _3476_/Y sky130_fd_sc_hd__nor2_1
X_5215_ _5369_/CLK _5215_/D vssd1 vssd1 vccd1 vccd1 _5215_/Q sky130_fd_sc_hd__dfxtp_1
X_5146_ _5313_/CLK _5146_/D vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5077_ _5077_/CLK _5077_/D vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dfxtp_1
X_4028_ _2833_/X _4022_/Y _2846_/X vssd1 vssd1 vccd1 vccd1 _4028_/X sky130_fd_sc_hd__o21a_1
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3330_ _4073_/D _3358_/A vssd1 vssd1 vccd1 vccd1 _3341_/B sky130_fd_sc_hd__nand2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _3305_/B _3261_/B vssd1 vssd1 vccd1 vccd1 _3309_/B sky130_fd_sc_hd__and2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5323_/CLK _5000_/D vssd1 vssd1 vccd1 vccd1 _5000_/Q sky130_fd_sc_hd__dfxtp_1
X_3192_ _3445_/C _3284_/A vssd1 vssd1 vccd1 vccd1 _3192_/Y sky130_fd_sc_hd__nand2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2976_ _5306_/Q _3075_/B _3074_/A vssd1 vssd1 vccd1 vccd1 _2976_/X sky130_fd_sc_hd__a21o_1
X_4715_ _4714_/A _4714_/B _5331_/Q vssd1 vssd1 vccd1 vccd1 _4716_/B sky130_fd_sc_hd__a21o_1
X_4646_ _5313_/Q _4644_/X _4662_/S vssd1 vssd1 vccd1 vccd1 _4647_/B sky130_fd_sc_hd__mux2_1
X_4577_ _5298_/Q _4577_/B vssd1 vssd1 vccd1 vccd1 _4577_/X sky130_fd_sc_hd__or2_1
X_3528_ _3528_/A _4730_/B vssd1 vssd1 vccd1 vccd1 _3658_/B sky130_fd_sc_hd__or2_1
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3459_ _3448_/Y _3456_/X _3458_/X vssd1 vssd1 vccd1 vccd1 _3459_/Y sky130_fd_sc_hd__a21oi_1
X_5129_ _5132_/CLK _5129_/D vssd1 vssd1 vccd1 vccd1 _5129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2830_ _5132_/Q _3462_/B _2859_/S vssd1 vssd1 vccd1 vccd1 _2830_/X sky130_fd_sc_hd__o21ba_1
XFILLER_43_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2761_ _4685_/A vssd1 vssd1 vccd1 vccd1 _2761_/X sky130_fd_sc_hd__clkbuf_2
X_2692_ _2695_/A vssd1 vssd1 vccd1 vccd1 _2692_/Y sky130_fd_sc_hd__inv_2
X_4500_ _4500_/A vssd1 vssd1 vccd1 vccd1 _5269_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA_1 _3431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4431_ _4165_/A _3659_/B _4429_/Y _4430_/Y _4093_/A vssd1 vssd1 vccd1 vccd1 _5245_/D
+ sky130_fd_sc_hd__a311o_1
X_4362_ _4402_/A vssd1 vssd1 vccd1 vccd1 _4362_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3313_ _3318_/A _3313_/B _3411_/B vssd1 vssd1 vccd1 vccd1 _3412_/B sky130_fd_sc_hd__and3b_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4293_ _4291_/X _5214_/Q _4309_/S vssd1 vssd1 vccd1 vccd1 _4294_/A sky130_fd_sc_hd__mux2_1
X_3244_ _5054_/Q _5053_/Q _3244_/C vssd1 vssd1 vccd1 vccd1 _3247_/C sky130_fd_sc_hd__or3_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _3074_/X _2889_/A _3076_/X _5317_/Q vssd1 vssd1 vccd1 vccd1 _3176_/B sky130_fd_sc_hd__a22o_1
XFILLER_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2959_ _5235_/Q vssd1 vssd1 vccd1 vccd1 _3090_/A sky130_fd_sc_hd__inv_2
XFILLER_136_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4629_ _4629_/A vssd1 vssd1 vccd1 vccd1 _5309_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4980_ _5453_/Q _4980_/B vssd1 vssd1 vccd1 vccd1 _4980_/X sky130_fd_sc_hd__or2_1
XFILLER_16_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3931_ _5085_/Q _3909_/X _3930_/X vssd1 vssd1 vccd1 vccd1 _5085_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3862_ hold40/A _2990_/X _5133_/D vssd1 vssd1 vccd1 vccd1 _3863_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5601_ _5601_/A _2633_/Y vssd1 vssd1 vccd1 vccd1 io_out[35] sky130_fd_sc_hd__ebufn_8
X_2813_ _2824_/S _2813_/B vssd1 vssd1 vccd1 vccd1 _2813_/Y sky130_fd_sc_hd__nor2_1
X_3793_ _5042_/Q _5041_/Q _5043_/Q vssd1 vssd1 vccd1 vccd1 _3794_/B sky130_fd_sc_hd__a21o_1
X_2744_ _4022_/A _2744_/B vssd1 vssd1 vccd1 vccd1 _2744_/X sky130_fd_sc_hd__and2_1
X_2675_ _2677_/A vssd1 vssd1 vccd1 vccd1 _2675_/Y sky130_fd_sc_hd__inv_2
X_5394_ _5403_/Q _5394_/D vssd1 vssd1 vccd1 vccd1 _5394_/Q sky130_fd_sc_hd__dfxtp_1
X_4414_ _5204_/Q _5174_/Q _4418_/S vssd1 vssd1 vccd1 vccd1 _4415_/B sky130_fd_sc_hd__mux2_1
X_4345_ _4345_/A vssd1 vssd1 vccd1 vccd1 _5225_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_59_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4276_ _4276_/A vssd1 vssd1 vccd1 vccd1 _4276_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3227_ _4990_/Q _4073_/B _3213_/Y vssd1 vssd1 vccd1 vccd1 _3238_/A sky130_fd_sc_hd__o21ba_2
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3158_ _3648_/A _3158_/B vssd1 vssd1 vccd1 vccd1 _3163_/A sky130_fd_sc_hd__xnor2_1
XFILLER_36_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ _5380_/Q _3028_/X _4833_/B _3009_/X _3088_/X vssd1 vssd1 vccd1 vccd1 _5380_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5504__94 vssd1 vssd1 vccd1 vccd1 _5504__94/HI _5607_/A sky130_fd_sc_hd__conb_1
XFILLER_58_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_11_wb_clk_i clkbuf_2_3_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5160_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4130_ _4130_/A vssd1 vssd1 vccd1 vccd1 _5166_/D sky130_fd_sc_hd__clkbuf_1
X_4061_ _5379_/Q hold61/A _4065_/S vssd1 vssd1 vccd1 vccd1 _4062_/A sky130_fd_sc_hd__mux2_1
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3012_ _5376_/Q _2925_/X _4832_/A _3009_/X _3011_/X vssd1 vssd1 vccd1 vccd1 _5376_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_36_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4963_ _4975_/A vssd1 vssd1 vccd1 vccd1 _4965_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3914_ _3919_/A vssd1 vssd1 vccd1 vccd1 _3915_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_32_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4894_ _4897_/B _4893_/Y _4841_/B vssd1 vssd1 vccd1 vccd1 _4894_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3845_ _3824_/C _3841_/X _3854_/A vssd1 vssd1 vccd1 vccd1 _3845_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_20_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3776_ _3729_/A _3776_/A2 _3764_/S _3192_/Y _3750_/X vssd1 vssd1 vccd1 vccd1 _3776_/X
+ sky130_fd_sc_hd__a32o_1
X_2727_ _2727_/A _4075_/A vssd1 vssd1 vccd1 vccd1 _2768_/B sky130_fd_sc_hd__nor2_1
X_5446_ _5446_/CLK _5446_/D vssd1 vssd1 vccd1 vccd1 _5446_/Q sky130_fd_sc_hd__dfxtp_1
X_2658_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2658_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5377_ _5403_/Q _5377_/D vssd1 vssd1 vccd1 vccd1 _5377_/Q sky130_fd_sc_hd__dfxtp_4
X_2589_ _2591_/A vssd1 vssd1 vccd1 vccd1 _2589_/Y sky130_fd_sc_hd__inv_2
X_4328_ _4328_/A _4328_/B vssd1 vssd1 vccd1 vccd1 _4681_/A sky130_fd_sc_hd__nor2_1
XFILLER_47_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4259_ _4609_/A _4259_/B vssd1 vssd1 vccd1 vccd1 _4260_/A sky130_fd_sc_hd__and2_1
XFILLER_28_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4006__1 _5132_/CLK vssd1 vssd1 vccd1 vccd1 _5120_/CLK sky130_fd_sc_hd__inv_2
XFILLER_7_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630_ _5001_/Q vssd1 vssd1 vccd1 vccd1 _3891_/B sky130_fd_sc_hd__clkbuf_2
X_3561_ _3563_/B _3563_/C _3569_/A vssd1 vssd1 vccd1 vccd1 _3561_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5300_ _5437_/CLK _5300_/D vssd1 vssd1 vccd1 vccd1 _5300_/Q sky130_fd_sc_hd__dfxtp_1
X_3492_ _4355_/C vssd1 vssd1 vccd1 vccd1 _4739_/A sky130_fd_sc_hd__buf_2
X_5231_ _5445_/CLK _5231_/D vssd1 vssd1 vccd1 vccd1 _5231_/Q sky130_fd_sc_hd__dfxtp_1
X_5162_ _5339_/CLK _5162_/D vssd1 vssd1 vccd1 vccd1 _5162_/Q sky130_fd_sc_hd__dfxtp_1
X_5093_ _5305_/CLK _5093_/D vssd1 vssd1 vccd1 vccd1 _5093_/Q sky130_fd_sc_hd__dfxtp_1
X_4113_ _5438_/Q _5336_/Q _5444_/Q vssd1 vssd1 vccd1 vccd1 _4113_/X sky130_fd_sc_hd__mux2_1
X_5495__85 vssd1 vssd1 vccd1 vccd1 _5495__85/HI _5573_/A sky130_fd_sc_hd__conb_1
X_4044_ _4044_/A vssd1 vssd1 vccd1 vccd1 _4071_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4946_ _4954_/A _4946_/B _4947_/B vssd1 vssd1 vccd1 vccd1 _5439_/D sky130_fd_sc_hd__nor3_1
X_4877_ _4880_/B _4876_/Y _4851_/X vssd1 vssd1 vccd1 vccd1 _4877_/Y sky130_fd_sc_hd__o21ai_1
X_3828_ _3828_/A _3828_/B vssd1 vssd1 vccd1 vccd1 _5052_/D sky130_fd_sc_hd__nor2_1
XFILLER_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3759_ _3751_/B _3758_/X _3277_/B vssd1 vssd1 vccd1 vccd1 _3759_/X sky130_fd_sc_hd__a21o_1
XFILLER_4_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5429_ _5430_/CLK _5429_/D vssd1 vssd1 vccd1 vccd1 _5429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4800_ _4800_/A vssd1 vssd1 vccd1 vccd1 _5390_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_15_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2992_ _2903_/B _2925_/X _2990_/X _2944_/X _2991_/X vssd1 vssd1 vccd1 vccd1 _5375_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _5370_/Q _5337_/Q vssd1 vssd1 vccd1 vccd1 _4731_/Y sky130_fd_sc_hd__nor2_1
X_4662_ _5317_/Q _4661_/X _4662_/S vssd1 vssd1 vccd1 vccd1 _4663_/B sky130_fd_sc_hd__mux2_1
X_3613_ _4587_/B _4328_/B vssd1 vssd1 vccd1 vccd1 _4504_/B sky130_fd_sc_hd__nor2_1
X_4593_ _5302_/Q _4081_/X _4586_/X _5324_/D vssd1 vssd1 vccd1 vccd1 _5302_/D sky130_fd_sc_hd__a22o_1
X_3544_ _5175_/Q _3541_/X _3543_/X _3535_/X vssd1 vssd1 vccd1 vccd1 _3545_/C sky130_fd_sc_hd__a22o_1
X_3475_ _3474_/X _5034_/Q _5033_/Q _5032_/Q _2795_/X _2846_/A vssd1 vssd1 vccd1 vccd1
+ _3475_/X sky130_fd_sc_hd__mux4_1
X_5214_ _5339_/CLK _5214_/D vssd1 vssd1 vccd1 vccd1 _5214_/Q sky130_fd_sc_hd__dfxtp_1
X_5145_ _5313_/CLK _5145_/D vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dfxtp_1
X_5076_ _5077_/CLK _5076_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4027_ _2833_/X _4022_/Y _4026_/Y vssd1 vssd1 vccd1 vccd1 _5127_/D sky130_fd_sc_hd__o21ai_1
XFILLER_44_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4929_ _4940_/S vssd1 vssd1 vccd1 vccd1 _4938_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_21_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _3260_/A _3551_/C _3260_/C _3260_/D vssd1 vssd1 vccd1 vccd1 _3261_/B sky130_fd_sc_hd__or4_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _3191_/A vssd1 vssd1 vccd1 vccd1 _3284_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5465__55 vssd1 vssd1 vccd1 vccd1 _5465__55/HI _5542_/A sky130_fd_sc_hd__conb_1
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2975_ _2975_/A vssd1 vssd1 vccd1 vccd1 _3074_/A sky130_fd_sc_hd__clkbuf_2
X_4714_ _4714_/A _4714_/B _5331_/Q vssd1 vssd1 vccd1 vccd1 _4722_/C sky130_fd_sc_hd__and3_1
X_4645_ _4666_/S vssd1 vssd1 vccd1 vccd1 _4662_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_30_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4576_ _5293_/Q _4566_/X _4575_/X _4571_/X vssd1 vssd1 vccd1 vccd1 _5297_/D sky130_fd_sc_hd__o211a_1
X_3527_ _4449_/C _4434_/B vssd1 vssd1 vccd1 vccd1 _3529_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3458_ _2846_/X _3462_/B _3457_/Y vssd1 vssd1 vccd1 vccd1 _3458_/X sky130_fd_sc_hd__o21a_1
X_3389_ _3369_/Y _3387_/X _3395_/A vssd1 vssd1 vccd1 vccd1 _3389_/Y sky130_fd_sc_hd__o21ai_1
X_5128_ _5132_/CLK _5128_/D vssd1 vssd1 vccd1 vccd1 _5128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5059_ _5439_/CLK _5059_/D vssd1 vssd1 vccd1 vccd1 _5059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2760_ _2760_/A _2768_/A _2760_/C vssd1 vssd1 vccd1 vccd1 _2760_/Y sky130_fd_sc_hd__nand3_1
X_2691_ _2695_/A vssd1 vssd1 vccd1 vccd1 _2691_/Y sky130_fd_sc_hd__inv_2
XANTENNA_2 _5639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4430_ _3659_/B _4429_/Y _5623_/A vssd1 vssd1 vccd1 vccd1 _4430_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_6_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4361_ _4739_/A _4363_/B _4363_/C vssd1 vssd1 vccd1 vccd1 _4402_/A sky130_fd_sc_hd__and3_1
X_3312_ _3308_/X _3356_/A _3355_/B vssd1 vssd1 vccd1 vccd1 _3388_/B sky130_fd_sc_hd__a21o_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4292_ _4292_/A vssd1 vssd1 vccd1 vccd1 _4309_/S sky130_fd_sc_hd__clkbuf_2
X_3243_ _3402_/A _3216_/A _3277_/B vssd1 vssd1 vccd1 vccd1 _3247_/B sky130_fd_sc_hd__a21oi_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _3648_/A _3174_/B vssd1 vssd1 vccd1 vccd1 _3179_/A sky130_fd_sc_hd__xnor2_1
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2958_ _2962_/A _2962_/B vssd1 vssd1 vccd1 vccd1 _2961_/B sky130_fd_sc_hd__xor2_1
XFILLER_136_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2889_ _2889_/A _2889_/B vssd1 vssd1 vccd1 vccd1 _2890_/A sky130_fd_sc_hd__nand2_1
X_4628_ _4632_/A _4628_/B vssd1 vssd1 vccd1 vccd1 _4629_/A sky130_fd_sc_hd__and2_1
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4559_ input3/X _4552_/X _4557_/X _4558_/X vssd1 vssd1 vccd1 vccd1 _5290_/D sky130_fd_sc_hd__o211a_1
XFILLER_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3930_ _5285_/Q _3910_/X _3697_/A _3929_/X vssd1 vssd1 vccd1 vccd1 _3930_/X sky130_fd_sc_hd__a211o_1
X_3861_ _3861_/A vssd1 vssd1 vccd1 vccd1 _5064_/D sky130_fd_sc_hd__clkbuf_1
X_5600_ _5600_/A _2632_/Y vssd1 vssd1 vccd1 vccd1 io_out[34] sky130_fd_sc_hd__ebufn_8
X_2812_ _2826_/A _2806_/X _2811_/X vssd1 vssd1 vccd1 vccd1 _2812_/Y sky130_fd_sc_hd__o21ai_1
X_3792_ _5042_/Q _5041_/Q _5043_/Q vssd1 vssd1 vccd1 vccd1 _3797_/B sky130_fd_sc_hd__and3_1
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2743_ _2743_/A _2752_/B _2752_/C vssd1 vssd1 vccd1 vccd1 _2744_/B sky130_fd_sc_hd__nor3_1
X_2674_ _2677_/A vssd1 vssd1 vccd1 vccd1 _2674_/Y sky130_fd_sc_hd__inv_2
X_5393_ _5403_/Q _5393_/D vssd1 vssd1 vccd1 vccd1 _5393_/Q sky130_fd_sc_hd__dfxtp_1
X_4413_ _3155_/B _4402_/X _4412_/X _4397_/X vssd1 vssd1 vccd1 vccd1 _5240_/D sky130_fd_sc_hd__o211a_1
X_4344_ _4348_/A _4344_/B vssd1 vssd1 vccd1 vccd1 _4345_/A sky130_fd_sc_hd__or2_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4275_ _4275_/A vssd1 vssd1 vccd1 vccd1 _4275_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _4991_/Q vssd1 vssd1 vccd1 vccd1 _4073_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3157_ _3647_/A _5400_/Q vssd1 vssd1 vccd1 vccd1 _3158_/B sky130_fd_sc_hd__and2_1
XFILLER_27_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3088_ _3106_/A _3652_/A vssd1 vssd1 vccd1 vccd1 _3088_/X sky130_fd_sc_hd__or2_1
XFILLER_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4060_ _4060_/A vssd1 vssd1 vccd1 vccd1 _5141_/D sky130_fd_sc_hd__clkbuf_1
X_3011_ _3106_/A _5232_/Q vssd1 vssd1 vccd1 vccd1 _3011_/X sky130_fd_sc_hd__or2_1
XFILLER_52_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4962_ _5243_/Q _5231_/Q vssd1 vssd1 vccd1 vccd1 _4975_/A sky130_fd_sc_hd__and2_1
X_4893_ _5416_/Q _4893_/B vssd1 vssd1 vccd1 vccd1 _4893_/Y sky130_fd_sc_hd__nor2_1
X_3913_ _3913_/A vssd1 vssd1 vccd1 vccd1 _3919_/A sky130_fd_sc_hd__clkbuf_2
X_3844_ _3844_/A vssd1 vssd1 vccd1 vccd1 _5057_/D sky130_fd_sc_hd__clkbuf_1
X_3775_ _5030_/Q _3767_/X _3740_/X _3774_/X vssd1 vssd1 vccd1 vccd1 _5030_/D sky130_fd_sc_hd__a22o_1
X_2726_ _3596_/A _3720_/B vssd1 vssd1 vccd1 vccd1 _4075_/A sky130_fd_sc_hd__or2_1
X_2657_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2657_/Y sky130_fd_sc_hd__inv_2
X_5445_ _5445_/CLK _5445_/D vssd1 vssd1 vccd1 vccd1 _5445_/Q sky130_fd_sc_hd__dfxtp_1
X_5376_ _5403_/Q _5376_/D vssd1 vssd1 vccd1 vccd1 _5376_/Q sky130_fd_sc_hd__dfxtp_4
X_2588_ _2591_/A vssd1 vssd1 vccd1 vccd1 _2588_/Y sky130_fd_sc_hd__inv_2
X_4327_ _4693_/B _4333_/B _3693_/B vssd1 vssd1 vccd1 vccd1 _4327_/X sky130_fd_sc_hd__a21o_1
X_4258_ _5206_/Q _5202_/Q _4258_/S vssd1 vssd1 vccd1 vccd1 _4259_/B sky130_fd_sc_hd__mux2_1
X_3209_ _4995_/Q _4996_/Q vssd1 vssd1 vccd1 vccd1 _3292_/A sky130_fd_sc_hd__or2_1
XFILLER_27_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4189_ _4189_/A vssd1 vssd1 vccd1 vccd1 _5185_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5531__121 vssd1 vssd1 vccd1 vccd1 _5531__121/HI _5531__121/LO sky130_fd_sc_hd__conb_1
XFILLER_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3560_ _3560_/A vssd1 vssd1 vccd1 vccd1 _4988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_5_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5230_ _5445_/CLK _5230_/D vssd1 vssd1 vccd1 vccd1 _5230_/Q sky130_fd_sc_hd__dfxtp_1
X_3491_ _5354_/Q vssd1 vssd1 vccd1 vccd1 _4355_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5161_ _5339_/CLK _5161_/D vssd1 vssd1 vccd1 vccd1 _5161_/Q sky130_fd_sc_hd__dfxtp_1
X_4112_ _4112_/A _4220_/C vssd1 vssd1 vccd1 vccd1 _4115_/B sky130_fd_sc_hd__nand2_2
X_5092_ _5322_/CLK _5092_/D vssd1 vssd1 vccd1 vccd1 _5092_/Q sky130_fd_sc_hd__dfxtp_1
X_4043_ _4043_/A _4043_/B vssd1 vssd1 vccd1 vccd1 _5132_/D sky130_fd_sc_hd__nor2_1
XFILLER_37_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4945_ _5444_/Q _5439_/Q _4945_/C vssd1 vssd1 vccd1 vccd1 _4947_/B sky130_fd_sc_hd__and3_1
XFILLER_33_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4876_ _5411_/Q _4875_/C _5412_/Q vssd1 vssd1 vccd1 vccd1 _4876_/Y sky130_fd_sc_hd__a21oi_1
X_3827_ _3829_/B _3829_/C _3826_/X vssd1 vssd1 vccd1 vccd1 _3828_/B sky130_fd_sc_hd__o21ai_1
X_3758_ _3841_/A _3847_/A vssd1 vssd1 vccd1 vccd1 _3758_/X sky130_fd_sc_hd__or2_1
X_2709_ _5118_/Q _5111_/Q vssd1 vssd1 vccd1 vccd1 _2729_/C sky130_fd_sc_hd__or2b_1
X_3689_ _5328_/Q _5327_/Q vssd1 vssd1 vccd1 vccd1 _4333_/B sky130_fd_sc_hd__or2_1
X_5428_ _5430_/CLK _5428_/D vssd1 vssd1 vccd1 vccd1 _5428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5359_ _5444_/CLK _5359_/D vssd1 vssd1 vccd1 vccd1 _5359_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5515__105 vssd1 vssd1 vccd1 vccd1 _5515__105/HI _5631_/A sky130_fd_sc_hd__conb_1
XFILLER_55_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2991_ _2991_/A _5231_/Q vssd1 vssd1 vccd1 vccd1 _2991_/X sky130_fd_sc_hd__or2_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _4730_/A _4730_/B vssd1 vssd1 vccd1 vccd1 _4942_/D sky130_fd_sc_hd__and2_1
X_4661_ _5299_/Q _5269_/Q _4661_/S vssd1 vssd1 vccd1 vccd1 _4661_/X sky130_fd_sc_hd__mux2_1
X_3612_ _5321_/Q vssd1 vssd1 vccd1 vccd1 _4328_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4592_ _4692_/C _4588_/X _4591_/Y _4350_/A vssd1 vssd1 vccd1 vccd1 _5324_/D sky130_fd_sc_hd__o211a_1
X_3543_ _5221_/Q _3543_/B vssd1 vssd1 vccd1 vccd1 _3543_/X sky130_fd_sc_hd__or2_1
X_3474_ _5031_/Q _3474_/B vssd1 vssd1 vccd1 vccd1 _3474_/X sky130_fd_sc_hd__and2_1
X_5213_ _5339_/CLK _5213_/D vssd1 vssd1 vccd1 vccd1 _5213_/Q sky130_fd_sc_hd__dfxtp_1
X_5144_ _5313_/CLK _5144_/D vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5075_ _5077_/CLK _5075_/D vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfxtp_1
X_4026_ _2833_/X _4022_/Y _4025_/Y vssd1 vssd1 vccd1 vccd1 _4026_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4928_ _4928_/A vssd1 vssd1 vccd1 vccd1 _5429_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_60_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4901_/A _4859_/B vssd1 vssd1 vccd1 vccd1 _4859_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _5060_/Q _5059_/Q _5058_/Q _5057_/Q _5061_/Q vssd1 vssd1 vccd1 vccd1 _3191_/A
+ sky130_fd_sc_hd__a41oi_4
XFILLER_54_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2974_ _2974_/A vssd1 vssd1 vccd1 vccd1 _3075_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_6_wb_clk_i clkbuf_2_1_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5443_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4713_ _4714_/A _4714_/B _4712_/Y vssd1 vssd1 vccd1 vccd1 _5330_/D sky130_fd_sc_hd__o21a_1
X_4644_ _5295_/Q _5265_/Q _4661_/S vssd1 vssd1 vccd1 vccd1 _4644_/X sky130_fd_sc_hd__mux2_1
X_4575_ _5297_/Q _4577_/B vssd1 vssd1 vccd1 vccd1 _4575_/X sky130_fd_sc_hd__or2_1
X_3526_ _3526_/A vssd1 vssd1 vccd1 vccd1 _4434_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3457_ _2846_/X _2822_/B _2838_/X vssd1 vssd1 vccd1 vccd1 _3457_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3388_ _3388_/A _3388_/B vssd1 vssd1 vccd1 vccd1 _3395_/A sky130_fd_sc_hd__xnor2_1
X_5127_ _5132_/CLK _5127_/D vssd1 vssd1 vccd1 vccd1 _5127_/Q sky130_fd_sc_hd__dfxtp_1
X_5058_ _5058_/CLK _5058_/D vssd1 vssd1 vccd1 vccd1 _5058_/Q sky130_fd_sc_hd__dfxtp_1
X_4009_ _5121_/Q vssd1 vssd1 vccd1 vccd1 _4012_/A sky130_fd_sc_hd__inv_2
XFILLER_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2690_ _2690_/A vssd1 vssd1 vccd1 vccd1 _2695_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_3 _5639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4360_ _4434_/A _4220_/C _4155_/X _3662_/X _3667_/A vssd1 vssd1 vccd1 vccd1 _4363_/C
+ sky130_fd_sc_hd__a32oi_4
X_3311_ _3354_/A _3354_/B vssd1 vssd1 vccd1 vccd1 _3355_/B sky130_fd_sc_hd__and2_1
XFILLER_6_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4291_ _5210_/Q _4275_/X _4290_/X vssd1 vssd1 vccd1 vccd1 _4291_/X sky130_fd_sc_hd__a21o_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3225_/X _3265_/B _3264_/A vssd1 vssd1 vccd1 vccd1 _3263_/A sky130_fd_sc_hd__a21oi_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3173_ _3647_/A _5401_/Q vssd1 vssd1 vccd1 vccd1 _3174_/B sky130_fd_sc_hd__and2_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2957_ _3033_/A _2957_/B vssd1 vssd1 vccd1 vccd1 _2962_/B sky130_fd_sc_hd__xnor2_1
X_2888_ _5240_/Q vssd1 vssd1 vccd1 vccd1 _2973_/A sky130_fd_sc_hd__clkbuf_2
X_4627_ _5309_/Q _4626_/X _4640_/S vssd1 vssd1 vccd1 vccd1 _4628_/B sky130_fd_sc_hd__mux2_1
X_4558_ _4571_/A vssd1 vssd1 vccd1 vccd1 _4558_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4489_ _4489_/A vssd1 vssd1 vccd1 vccd1 _5264_/D sky130_fd_sc_hd__clkbuf_1
X_3509_ _5253_/Q _5252_/Q vssd1 vssd1 vccd1 vccd1 _3510_/C sky130_fd_sc_hd__nor2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3860_ _5064_/Q _2965_/X _5133_/D vssd1 vssd1 vccd1 vccd1 _3861_/A sky130_fd_sc_hd__mux2_1
XFILLER_32_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2811_ _3464_/A _3461_/A _2810_/X vssd1 vssd1 vccd1 vccd1 _2811_/X sky130_fd_sc_hd__a21o_1
X_3791_ _3791_/A vssd1 vssd1 vccd1 vccd1 _5042_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_32_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2742_ _2753_/A vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2673_ _2677_/A vssd1 vssd1 vccd1 vccd1 _2673_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4412_ _4419_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4412_/X sky130_fd_sc_hd__or2_1
X_5392_ _5403_/Q _5392_/D vssd1 vssd1 vccd1 vccd1 _5392_/Q sky130_fd_sc_hd__dfxtp_1
X_4343_ _5578_/A _4342_/X _4347_/S vssd1 vssd1 vccd1 vccd1 _4344_/B sky130_fd_sc_hd__mux2_1
X_4274_ _4274_/A vssd1 vssd1 vccd1 vccd1 _5210_/D sky130_fd_sc_hd__clkbuf_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3225_ _3192_/Y _3224_/A _3215_/X _3224_/Y vssd1 vssd1 vccd1 vccd1 _3225_/X sky130_fd_sc_hd__a211o_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3156_ _5384_/Q _3028_/A _4834_/C _3120_/X _3155_/X vssd1 vssd1 vccd1 vccd1 _5384_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_36_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3087_ _3142_/A vssd1 vssd1 vccd1 vccd1 _3652_/A sky130_fd_sc_hd__buf_2
XFILLER_54_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3989_ _5108_/Q _3983_/A _3980_/A _4837_/B vssd1 vssd1 vccd1 vccd1 _5108_/D sky130_fd_sc_hd__a22o_1
XFILLER_58_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_wb_clk_i clkbuf_2_2_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5430_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_3_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3010_ _4791_/A vssd1 vssd1 vccd1 vccd1 _3106_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_37_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4961_ _5446_/Q _4959_/X _2787_/B vssd1 vssd1 vccd1 vccd1 _5446_/D sky130_fd_sc_hd__a21o_1
X_4892_ _5416_/Q _4893_/B vssd1 vssd1 vccd1 vccd1 _4897_/B sky130_fd_sc_hd__and2_1
X_3912_ _3912_/A _3912_/B vssd1 vssd1 vccd1 vccd1 _3913_/A sky130_fd_sc_hd__nor2_1
X_3843_ _3841_/X _3854_/A _3843_/C vssd1 vssd1 vccd1 vccd1 _3844_/A sky130_fd_sc_hd__and3b_1
XFILLER_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3774_ _3741_/X _3772_/Y _3773_/X _3606_/A vssd1 vssd1 vccd1 vccd1 _3774_/X sky130_fd_sc_hd__a22o_1
XFILLER_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2725_ _2753_/A _2725_/B vssd1 vssd1 vccd1 vccd1 _3720_/B sky130_fd_sc_hd__or2_2
X_5444_ _5444_/CLK _5444_/D vssd1 vssd1 vccd1 vccd1 _5444_/Q sky130_fd_sc_hd__dfxtp_2
X_2656_ _2659_/A vssd1 vssd1 vccd1 vccd1 _2656_/Y sky130_fd_sc_hd__inv_2
X_5375_ _5403_/Q _5375_/D vssd1 vssd1 vccd1 vccd1 _5375_/Q sky130_fd_sc_hd__dfxtp_1
X_2587_ _2591_/A vssd1 vssd1 vccd1 vccd1 _2587_/Y sky130_fd_sc_hd__inv_2
X_4326_ _4589_/A vssd1 vssd1 vccd1 vccd1 _4693_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4257_ _4257_/A vssd1 vssd1 vccd1 vccd1 _5205_/D sky130_fd_sc_hd__clkbuf_1
X_3208_ _4992_/Q _4993_/Q _4994_/Q vssd1 vssd1 vccd1 vccd1 _3211_/A sky130_fd_sc_hd__o21a_1
X_4188_ _4187_/X _5185_/Q _4197_/S vssd1 vssd1 vccd1 vccd1 _4189_/A sky130_fd_sc_hd__mux2_1
X_3139_ _3139_/A _3139_/B vssd1 vssd1 vccd1 vccd1 _3148_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_136_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3490_ _3490_/A vssd1 vssd1 vccd1 vccd1 _5591_/A sky130_fd_sc_hd__clkbuf_1
X_5160_ _5160_/CLK _5160_/D vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4111_ hold37/A _4109_/A _4110_/Y vssd1 vssd1 vccd1 vccd1 _5160_/D sky130_fd_sc_hd__o21a_1
X_5091_ _5322_/CLK _5091_/D vssd1 vssd1 vccd1 vccd1 _5091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4042_ _4042_/A _4042_/B vssd1 vssd1 vccd1 vccd1 _4043_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4944_ _4789_/A _4945_/C _5439_/Q vssd1 vssd1 vccd1 vccd1 _4946_/B sky130_fd_sc_hd__a21oi_1
XFILLER_40_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4875_ _5411_/Q _5412_/Q _4875_/C vssd1 vssd1 vccd1 vccd1 _4880_/B sky130_fd_sc_hd__and3_1
XFILLER_137_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3826_ _3838_/A vssd1 vssd1 vccd1 vccd1 _3826_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3757_ _3757_/A vssd1 vssd1 vccd1 vccd1 _5026_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2708_ _5113_/Q _5112_/Q _2752_/B vssd1 vssd1 vccd1 vccd1 _3705_/D sky130_fd_sc_hd__or3_1
X_3688_ _5325_/Q vssd1 vssd1 vccd1 vccd1 _4692_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_2639_ _2640_/A vssd1 vssd1 vccd1 vccd1 _2639_/Y sky130_fd_sc_hd__inv_2
X_5427_ _5430_/CLK _5427_/D vssd1 vssd1 vccd1 vccd1 _5427_/Q sky130_fd_sc_hd__dfxtp_1
X_5358_ _5444_/CLK _5358_/D vssd1 vssd1 vccd1 vccd1 _5358_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4309_ _4308_/X _5218_/Q _4309_/S vssd1 vssd1 vccd1 vccd1 _4310_/A sky130_fd_sc_hd__mux2_1
X_5486__76 vssd1 vssd1 vccd1 vccd1 _5486__76/HI _5564_/A sky130_fd_sc_hd__conb_1
XFILLER_28_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5289_ _5437_/CLK _5289_/D vssd1 vssd1 vccd1 vccd1 _5289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_137_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2990_ _4831_/D vssd1 vssd1 vccd1 vccd1 _2990_/X sky130_fd_sc_hd__clkbuf_4
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4660_ _4660_/A vssd1 vssd1 vccd1 vccd1 _5316_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_30_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3611_ _5322_/Q vssd1 vssd1 vccd1 vccd1 _4587_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_4591_ _4591_/A _4591_/B vssd1 vssd1 vccd1 vccd1 _4591_/Y sky130_fd_sc_hd__nand2_1
X_3542_ _3547_/B vssd1 vssd1 vccd1 vccd1 _3543_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3473_ _3465_/Y _3469_/X _3470_/Y _4038_/B vssd1 vssd1 vccd1 vccd1 _3473_/Y sky130_fd_sc_hd__o211ai_1
X_5212_ _5339_/CLK _5212_/D vssd1 vssd1 vccd1 vccd1 _5212_/Q sky130_fd_sc_hd__dfxtp_1
X_5143_ _5313_/CLK _5143_/D vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5074_ _5077_/CLK _5074_/D vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4025_ _4033_/A vssd1 vssd1 vccd1 vccd1 _4025_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4927_ _5429_/Q _5380_/Q _4927_/S vssd1 vssd1 vccd1 vccd1 _4928_/A sky130_fd_sc_hd__mux2_1
XFILLER_33_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4858_ _5408_/Q _4864_/C vssd1 vssd1 vccd1 vccd1 _4859_/B sky130_fd_sc_hd__xnor2_1
X_3809_ _3809_/A _3809_/B vssd1 vssd1 vccd1 vccd1 _5047_/D sky130_fd_sc_hd__nor2_1
X_4789_ _4789_/A _4789_/B _4789_/C vssd1 vssd1 vccd1 vccd1 _4790_/A sky130_fd_sc_hd__and3_1
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_137_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2973_ _2973_/A vssd1 vssd1 vccd1 vccd1 _3155_/B sky130_fd_sc_hd__clkbuf_2
X_4712_ _4714_/A _4714_/B _4710_/B vssd1 vssd1 vccd1 vccd1 _4712_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_30_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4643_ _4665_/S vssd1 vssd1 vccd1 vccd1 _4661_/S sky130_fd_sc_hd__clkbuf_2
X_4574_ _5292_/Q _4566_/X _4573_/X _4571_/X vssd1 vssd1 vccd1 vccd1 _5296_/D sky130_fd_sc_hd__o211a_1
X_3525_ _5249_/Q vssd1 vssd1 vccd1 vccd1 _4449_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_3456_ _2859_/X _2855_/X _2856_/X _2858_/X _2846_/X _4034_/A vssd1 vssd1 vccd1 vccd1
+ _3456_/X sky130_fd_sc_hd__mux4_1
X_3387_ _3393_/B _3387_/B _3387_/C vssd1 vssd1 vccd1 vccd1 _3387_/X sky130_fd_sc_hd__and3_1
X_5126_ _5126_/CLK _5126_/D vssd1 vssd1 vccd1 vccd1 _5126_/Q sky130_fd_sc_hd__dfxtp_1
X_5057_ _5058_/CLK _5057_/D vssd1 vssd1 vccd1 vccd1 _5057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4008_ _4024_/A vssd1 vssd1 vccd1 vccd1 _5122_/D sky130_fd_sc_hd__clkinv_2
XFILLER_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_136_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_44_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5470__60 vssd1 vssd1 vccd1 vccd1 _5470__60/HI _5547_/A sky130_fd_sc_hd__conb_1
XFILLER_16_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_4 _5640_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_137_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3310_ _3263_/A _3263_/B _3309_/Y vssd1 vssd1 vccd1 vccd1 _3356_/A sky130_fd_sc_hd__o21ai_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4290_ _5164_/Q _4285_/X _4276_/X _5190_/Q vssd1 vssd1 vccd1 vccd1 _4290_/X sky130_fd_sc_hd__a22o_1
X_3241_ _3192_/Y _3252_/S _3215_/X _3240_/Y vssd1 vssd1 vccd1 vccd1 _3264_/A sky130_fd_sc_hd__o211a_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3172_ _2889_/B _3028_/A _3170_/X _3120_/X _3171_/X vssd1 vssd1 vccd1 vccd1 _5385_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_19_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2956_ _2973_/A _2903_/C _2955_/X _2980_/A vssd1 vssd1 vccd1 vccd1 _2957_/B sky130_fd_sc_hd__o211a_1
X_2887_ _5236_/Q vssd1 vssd1 vccd1 vccd1 _3033_/A sky130_fd_sc_hd__buf_2
X_4626_ _5291_/Q _5261_/Q _4639_/S vssd1 vssd1 vccd1 vccd1 _4626_/X sky130_fd_sc_hd__mux2_1
X_4557_ _5290_/Q _4564_/B vssd1 vssd1 vccd1 vccd1 _4557_/X sky130_fd_sc_hd__or2_1
X_3508_ _5250_/Q vssd1 vssd1 vccd1 vccd1 _3510_/B sky130_fd_sc_hd__clkinv_2
X_4488_ _5264_/Q _5102_/Q _4492_/S vssd1 vssd1 vccd1 vccd1 _4489_/A sky130_fd_sc_hd__mux2_1
X_3439_ _4073_/C _4074_/B _3578_/B _3439_/D vssd1 vssd1 vccd1 vccd1 _3440_/A sky130_fd_sc_hd__or4_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5446_/CLK _5109_/D vssd1 vssd1 vccd1 vccd1 _5109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2810_ _5029_/Q _5030_/Q _2872_/S vssd1 vssd1 vccd1 vccd1 _2810_/X sky130_fd_sc_hd__mux2_1
X_3790_ _2518_/Y _3820_/A vssd1 vssd1 vccd1 vccd1 _3791_/A sky130_fd_sc_hd__and2b_1
X_2741_ _3754_/A vssd1 vssd1 vccd1 vccd1 _3729_/A sky130_fd_sc_hd__clkbuf_2
X_2672_ _2690_/A vssd1 vssd1 vccd1 vccd1 _2677_/A sky130_fd_sc_hd__buf_2
X_4411_ _5203_/Q _5173_/Q _4418_/S vssd1 vssd1 vccd1 vccd1 _4412_/B sky130_fd_sc_hd__mux2_1
X_5391_ _5403_/Q _5391_/D vssd1 vssd1 vccd1 vccd1 _5391_/Q sky130_fd_sc_hd__dfxtp_1
X_4342_ _5269_/Q _3919_/A _3943_/X _5091_/Q _3947_/A vssd1 vssd1 vccd1 vccd1 _4342_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_59_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4273_ _4272_/X _5210_/Q _4288_/S vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__mux2_1
X_3224_ _3224_/A _3240_/B vssd1 vssd1 vccd1 vccd1 _3224_/Y sky130_fd_sc_hd__nor2_1
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

